//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  AND3_X1   g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT66), .Z(new_n214));
  AOI21_X1  g0014(.A(new_n207), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT67), .Z(new_n218));
  INV_X1    g0018(.A(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n207), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n222), .A2(new_n223), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n229), .B1(new_n223), .B2(new_n222), .C1(new_n216), .C2(new_n215), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n218), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n251), .B1(new_n254), .B2(G226), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT69), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1698), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT70), .B(G223), .Z(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n260), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n267), .A2(G222), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n252), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n256), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n224), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n225), .A2(G33), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n276), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n219), .A2(new_n225), .A3(G1), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n275), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G1), .B2(new_n225), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G50), .ZN(new_n286));
  INV_X1    g0086(.A(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n202), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n282), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n270), .A2(G169), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n273), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT72), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n251), .B1(new_n254), .B2(G238), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n267), .A2(G226), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n266), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G232), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G97), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n293), .B1(new_n299), .B2(new_n253), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(KEYINPUT75), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(KEYINPUT75), .B2(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G169), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n307));
  NAND2_X1  g0107(.A1(KEYINPUT76), .A2(KEYINPUT13), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n300), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G179), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n264), .B2(new_n278), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n312), .B2(new_n285), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT11), .B1(new_n314), .B2(new_n275), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n219), .A2(G1), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(G20), .A3(new_n312), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT12), .Z(new_n320));
  NOR3_X1   g0120(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n304), .A2(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n309), .A2(G190), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n312), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n201), .ZN(new_n330));
  INV_X1    g0130(.A(G159), .ZN(new_n331));
  INV_X1    g0131(.A(new_n280), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n261), .B2(G20), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n312), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n333), .B1(new_n337), .B2(KEYINPUT77), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(KEYINPUT77), .B2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT16), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n258), .A2(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n260), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n258), .A2(KEYINPUT78), .ZN(new_n344));
  OAI211_X1 g0144(.A(KEYINPUT7), .B(new_n225), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n312), .B1(new_n345), .B2(new_n335), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n340), .B1(new_n346), .B2(new_n333), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n275), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n284), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n277), .B1(new_n248), .B2(G20), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(KEYINPUT79), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(KEYINPUT79), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n351), .A2(new_n352), .B1(new_n283), .B2(new_n277), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n251), .B1(new_n254), .B2(G232), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n296), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n267), .A2(G223), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n354), .B1(new_n357), .B2(new_n253), .ZN(new_n358));
  INV_X1    g0158(.A(G200), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G190), .B2(new_n358), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n348), .A2(new_n353), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT17), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n348), .A2(new_n353), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n358), .A2(G179), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n358), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT18), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n362), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n364), .A2(new_n370), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n270), .A2(G190), .ZN(new_n376));
  XOR2_X1   g0176(.A(new_n289), .B(KEYINPUT9), .Z(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(new_n359), .C2(new_n270), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT10), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n267), .A2(G232), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT73), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n296), .A2(G238), .B1(G107), .B2(new_n266), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n253), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n254), .A2(G244), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n250), .B2(new_n249), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G200), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n283), .A2(G77), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n285), .B2(G77), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n392), .A2(new_n278), .B1(new_n225), .B2(new_n264), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n277), .B(KEYINPUT74), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(new_n280), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n391), .B1(new_n397), .B2(new_n275), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n386), .A2(G179), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n383), .B2(new_n385), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n379), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n292), .A2(new_n327), .A3(new_n375), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n258), .A2(new_n260), .A3(G244), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(G1698), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(new_n258), .A3(new_n260), .A4(G244), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G283), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n258), .A2(new_n260), .A3(G250), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n295), .B1(new_n414), .B2(KEYINPUT4), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT80), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(KEYINPUT4), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT80), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n407), .A2(new_n408), .B1(G33), .B2(G283), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n411), .A4(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n252), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G41), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT81), .B1(new_n423), .B2(KEYINPUT5), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT5), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(G41), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n248), .A2(G45), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n425), .A2(G41), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(KEYINPUT81), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n252), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G257), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n429), .A3(G274), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n422), .A2(G179), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n422), .A2(new_n433), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n367), .ZN(new_n436));
  INV_X1    g0236(.A(G107), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n345), .B2(new_n335), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT6), .ZN(new_n439));
  INV_X1    g0239(.A(G97), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n437), .ZN(new_n441));
  NOR2_X1   g0241(.A1(G97), .A2(G107), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n437), .A2(KEYINPUT6), .A3(G97), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n445), .A2(new_n225), .B1(new_n264), .B2(new_n332), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n275), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n287), .A2(G97), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n284), .B1(G1), .B2(new_n257), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT82), .B1(new_n436), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n422), .A2(G179), .A3(new_n433), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n367), .B1(new_n422), .B2(new_n433), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(KEYINPUT82), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n452), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n435), .A2(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n422), .A2(new_n433), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G190), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n296), .A2(G264), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n261), .A2(G257), .A3(new_n295), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n266), .A2(G303), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n253), .B1(new_n470), .B2(KEYINPUT85), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n430), .A2(G270), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n432), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT84), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n478), .A3(new_n432), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n257), .A2(G97), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(new_n482), .B2(new_n412), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n225), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n275), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g0286(.A(new_n486), .B(KEYINPUT20), .Z(new_n487));
  NAND2_X1  g0287(.A1(new_n287), .A2(new_n484), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n450), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n481), .A2(KEYINPUT21), .A3(G169), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n471), .A2(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(G169), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(G179), .A3(new_n490), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n481), .A2(new_n359), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n387), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n392), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n287), .ZN(new_n503));
  NAND3_X1  g0303(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n504), .A2(new_n505), .A3(new_n225), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n504), .B2(new_n225), .ZN(new_n507));
  INV_X1    g0307(.A(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n440), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n506), .A2(new_n507), .B1(G107), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n261), .A2(new_n225), .A3(G68), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n298), .A2(G20), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n511), .C1(KEYINPUT19), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n503), .B1(new_n513), .B2(new_n275), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n450), .A2(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n261), .A2(G238), .A3(new_n295), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n258), .A2(new_n260), .A3(G244), .A4(G1698), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n252), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n427), .A2(G250), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n248), .A2(G45), .A3(G274), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n252), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n359), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n520), .B2(new_n252), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n387), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n516), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n514), .B1(new_n392), .B2(new_n449), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n521), .A2(G179), .A3(new_n525), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n367), .B2(new_n528), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n535));
  INV_X1    g0335(.A(G294), .ZN(new_n536));
  OAI221_X1 g0336(.A(new_n535), .B1(new_n257), .B2(new_n536), .C1(G1698), .C2(new_n414), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n252), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n430), .A2(G264), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n432), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G169), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n271), .B2(new_n540), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n437), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT23), .B1(new_n437), .B2(G20), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n543), .A2(new_n544), .B1(G20), .B2(new_n518), .ZN(new_n545));
  OR4_X1    g0345(.A1(KEYINPUT22), .A2(new_n266), .A3(G20), .A4(new_n508), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n261), .A2(new_n225), .A3(G87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n276), .B1(new_n549), .B2(KEYINPUT24), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(KEYINPUT24), .B2(new_n549), .ZN(new_n551));
  INV_X1    g0351(.A(new_n318), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n437), .A2(G20), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT25), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OR3_X1    g0354(.A1(new_n552), .A2(KEYINPUT25), .A3(new_n553), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n449), .C2(new_n437), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n556), .B(KEYINPUT86), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n542), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n540), .A2(new_n359), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n540), .A2(G190), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n557), .B(new_n551), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n534), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n465), .A2(new_n501), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n406), .A2(new_n564), .ZN(G372));
  NAND2_X1  g0365(.A1(new_n370), .A2(new_n372), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n311), .A2(new_n322), .B1(new_n326), .B2(new_n402), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n364), .A2(new_n374), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n292), .B1(new_n570), .B2(new_n379), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT87), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n532), .B(new_n572), .C1(new_n367), .C2(new_n528), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n573), .A2(new_n531), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n528), .A2(new_n367), .ZN(new_n575));
  AOI211_X1 g0375(.A(new_n271), .B(new_n524), .C1(new_n520), .C2(new_n252), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT87), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n530), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n559), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n562), .B(new_n578), .C1(new_n497), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n464), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT88), .B1(new_n436), .B2(new_n452), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n452), .B(KEYINPUT88), .C1(new_n454), .C2(new_n455), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n578), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT26), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n527), .A2(new_n529), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n514), .A3(new_n515), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n533), .A2(new_n531), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n456), .ZN(new_n594));
  XOR2_X1   g0394(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n585), .A2(new_n586), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n577), .A2(new_n531), .A3(new_n573), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT90), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n534), .B(new_n596), .C1(new_n453), .C2(new_n457), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n588), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT88), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n591), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n604), .B2(new_n583), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n605), .B2(KEYINPUT26), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT90), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n598), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n581), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n571), .B1(new_n406), .B2(new_n609), .ZN(G369));
  OR3_X1    g0410(.A1(new_n552), .A2(KEYINPUT27), .A3(G20), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT27), .B1(new_n552), .B2(G20), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(G213), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G343), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n551), .B2(new_n557), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT91), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n562), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n559), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n579), .A2(new_n616), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n497), .A2(new_n616), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n579), .B2(new_n616), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n490), .A2(new_n615), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n497), .B2(new_n500), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n497), .B2(new_n628), .ZN(new_n630));
  INV_X1    g0430(.A(G330), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n624), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n627), .A2(new_n634), .ZN(G399));
  NAND2_X1  g0435(.A1(new_n221), .A2(new_n423), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n509), .A2(G107), .A3(G116), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G1), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n227), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT28), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n528), .A2(G179), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n481), .A2(new_n461), .A3(new_n540), .A4(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n576), .A2(new_n539), .A3(new_n538), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n493), .A2(new_n643), .A3(new_n435), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT30), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT92), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n647), .A4(new_n642), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n616), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n465), .A2(new_n501), .A3(new_n563), .A4(new_n616), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(KEYINPUT31), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n646), .A2(new_n648), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT31), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n657), .A3(new_n616), .ZN(new_n658));
  OAI21_X1  g0458(.A(G330), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n609), .A2(new_n615), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT29), .ZN(new_n662));
  INV_X1    g0462(.A(new_n581), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n585), .A2(new_n586), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n594), .A2(new_n596), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n598), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(KEYINPUT93), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n668));
  OAI211_X1 g0468(.A(KEYINPUT29), .B(new_n616), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n660), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n640), .B1(new_n670), .B2(G1), .ZN(G364));
  NOR2_X1   g0471(.A1(new_n219), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G45), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n636), .A2(G1), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n224), .B1(G20), .B2(new_n367), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n271), .A2(new_n359), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT98), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n225), .A2(G190), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G159), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT99), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT32), .ZN(new_n685));
  NAND2_X1  g0485(.A1(G20), .A2(G179), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT96), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n387), .A2(new_n359), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n387), .A2(G200), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI22_X1  g0493(.A1(G50), .A2(new_n690), .B1(new_n693), .B2(G58), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n387), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G200), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n694), .B1(new_n264), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT97), .Z(new_n699));
  NAND3_X1  g0499(.A1(new_n680), .A2(new_n271), .A3(G200), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n225), .A2(new_n387), .A3(new_n359), .A4(G179), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI221_X1 g0502(.A(new_n261), .B1(new_n437), .B2(new_n700), .C1(new_n702), .C2(new_n508), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n225), .B1(new_n679), .B2(G190), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n440), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n695), .A2(new_n359), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n703), .B(new_n705), .C1(G68), .C2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n685), .A2(new_n699), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(KEYINPUT100), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT100), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n701), .B(KEYINPUT101), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n682), .A2(G329), .B1(G303), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G326), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n689), .ZN(new_n715));
  INV_X1    g0515(.A(G283), .ZN(new_n716));
  INV_X1    g0516(.A(G322), .ZN(new_n717));
  OAI221_X1 g0517(.A(new_n266), .B1(new_n716), .B2(new_n700), .C1(new_n692), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(G311), .B2(new_n696), .ZN(new_n719));
  INV_X1    g0519(.A(new_n704), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G294), .ZN(new_n721));
  XNOR2_X1  g0521(.A(KEYINPUT33), .B(G317), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n706), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n708), .A2(new_n711), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n676), .B1(new_n710), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n676), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n221), .A2(G116), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n221), .A2(new_n266), .ZN(new_n733));
  INV_X1    g0533(.A(G45), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n242), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT94), .Z(new_n736));
  AOI211_X1 g0536(.A(new_n733), .B(new_n736), .C1(new_n734), .C2(new_n228), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n220), .A2(new_n266), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n732), .B(new_n737), .C1(G355), .C2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n726), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n630), .A2(new_n729), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n675), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n630), .A2(new_n631), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n674), .B1(new_n743), .B2(new_n632), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT102), .ZN(G396));
  NOR2_X1   g0546(.A1(new_n676), .A2(new_n727), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n674), .B1(new_n264), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n676), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n712), .A2(G107), .B1(G303), .B2(new_n690), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n536), .B2(new_n692), .ZN(new_n751));
  INV_X1    g0551(.A(new_n706), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n484), .A2(new_n697), .B1(new_n752), .B2(new_n716), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n266), .B1(new_n508), .B2(new_n700), .C1(new_n681), .C2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n751), .A2(new_n753), .A3(new_n755), .A4(new_n705), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n704), .A2(new_n328), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n700), .A2(new_n312), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n266), .B(new_n758), .C1(new_n712), .C2(G50), .ZN(new_n759));
  INV_X1    g0559(.A(G132), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n760), .B2(new_n681), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G137), .A2(new_n690), .B1(new_n693), .B2(G143), .ZN(new_n762));
  INV_X1    g0562(.A(G150), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n762), .B1(new_n697), .B2(new_n331), .C1(new_n763), .C2(new_n752), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT34), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n757), .B(new_n761), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n756), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n402), .A2(new_n616), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n398), .A2(new_n616), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n389), .B2(new_n398), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n769), .B1(new_n771), .B2(new_n402), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n748), .B1(new_n749), .B2(new_n768), .C1(new_n773), .C2(new_n728), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n661), .B(new_n773), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n659), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n674), .B1(new_n775), .B2(new_n659), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(G384));
  NAND2_X1  g0579(.A1(new_n339), .A2(new_n340), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n341), .A2(new_n275), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n613), .B1(new_n781), .B2(new_n353), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n375), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n613), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n368), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n353), .B2(new_n781), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT37), .B1(new_n786), .B2(new_n363), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n365), .A2(new_n784), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n369), .A2(new_n788), .A3(new_n362), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(KEYINPUT37), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n783), .A2(KEYINPUT38), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT38), .B1(new_n783), .B2(new_n790), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n323), .B(new_n326), .C1(new_n321), .C2(new_n616), .ZN(new_n795));
  INV_X1    g0595(.A(new_n326), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n322), .B(new_n615), .C1(new_n311), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n585), .A2(new_n586), .ZN(new_n799));
  AOI211_X1 g0599(.A(KEYINPUT90), .B(new_n599), .C1(new_n799), .C2(new_n601), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n607), .B1(new_n606), .B2(new_n598), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n663), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(new_n616), .A3(new_n773), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT104), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n803), .A2(new_n804), .A3(new_n769), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n803), .B2(new_n769), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT105), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n609), .A2(new_n615), .A3(new_n772), .ZN(new_n809));
  INV_X1    g0609(.A(new_n769), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT104), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n803), .A2(new_n804), .A3(new_n769), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT105), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n813), .A2(new_n814), .A3(new_n798), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n794), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT39), .B1(new_n792), .B2(new_n793), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n791), .A2(KEYINPUT106), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT106), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n783), .A2(new_n790), .A3(new_n819), .A4(KEYINPUT38), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n789), .B(KEYINPUT37), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n375), .A2(new_n365), .A3(new_n784), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n818), .B(new_n820), .C1(KEYINPUT38), .C2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n817), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n323), .A2(new_n615), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(new_n826), .B1(new_n566), .B2(new_n613), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n816), .A2(new_n828), .A3(KEYINPUT107), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT107), .ZN(new_n830));
  INV_X1    g0630(.A(new_n794), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n814), .B1(new_n813), .B2(new_n798), .ZN(new_n832));
  INV_X1    g0632(.A(new_n798), .ZN(new_n833));
  AOI211_X1 g0633(.A(KEYINPUT105), .B(new_n833), .C1(new_n811), .C2(new_n812), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n830), .B1(new_n835), .B2(new_n827), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n662), .A2(new_n405), .A3(new_n669), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n571), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n837), .B(new_n839), .Z(new_n840));
  INV_X1    g0640(.A(KEYINPUT40), .ZN(new_n841));
  INV_X1    g0641(.A(new_n655), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n653), .A2(KEYINPUT31), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n772), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n798), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n845), .B2(new_n794), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n824), .A2(KEYINPUT40), .A3(new_n798), .A4(new_n844), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n842), .A2(new_n843), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n405), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n848), .B(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n631), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n840), .A2(new_n852), .B1(new_n248), .B2(new_n672), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n840), .B2(new_n852), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n228), .B(G77), .C1(new_n328), .C2(new_n312), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n202), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n248), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n445), .ZN(new_n858));
  OAI211_X1 g0658(.A(G116), .B(new_n226), .C1(new_n858), .C2(KEYINPUT35), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(KEYINPUT35), .B2(new_n858), .ZN(new_n860));
  XNOR2_X1  g0660(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OR3_X1    g0662(.A1(new_n854), .A2(new_n857), .A3(new_n862), .ZN(G367));
  NOR2_X1   g0663(.A1(new_n733), .A2(new_n238), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n730), .B1(new_n221), .B2(new_n392), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n675), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n712), .A2(KEYINPUT46), .A3(G116), .ZN(new_n867));
  INV_X1    g0667(.A(new_n700), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n261), .B1(new_n868), .B2(G97), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n702), .A2(new_n484), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n867), .B(new_n869), .C1(KEYINPUT46), .C2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n720), .A2(G107), .B1(G294), .B2(new_n706), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n716), .B2(new_n697), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n871), .B(new_n873), .C1(G317), .C2(new_n682), .ZN(new_n874));
  INV_X1    g0674(.A(G303), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n875), .A2(new_n692), .B1(new_n689), .B2(new_n754), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT110), .Z(new_n877));
  NOR2_X1   g0677(.A1(new_n704), .A2(new_n312), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n682), .A2(G137), .B1(G58), .B2(new_n701), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n202), .B2(new_n697), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n878), .B(new_n880), .C1(G159), .C2(new_n706), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n692), .A2(new_n763), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n261), .B1(new_n700), .B2(new_n264), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT111), .Z(new_n884));
  AOI211_X1 g0684(.A(new_n882), .B(new_n884), .C1(G143), .C2(new_n690), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n874), .A2(new_n877), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n886), .A2(KEYINPUT47), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n749), .B1(new_n886), .B2(KEYINPUT47), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n866), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n516), .A2(new_n615), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n578), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT108), .ZN(new_n892));
  OR3_X1    g0692(.A1(new_n598), .A2(new_n892), .A3(new_n890), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n598), .B2(new_n890), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n729), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n465), .B1(new_n459), .B2(new_n616), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n436), .A2(new_n452), .A3(new_n615), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n626), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT42), .Z(new_n902));
  INV_X1    g0702(.A(new_n900), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n458), .B1(new_n903), .B2(new_n559), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n616), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n902), .A2(new_n905), .B1(KEYINPUT43), .B2(new_n895), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n903), .A2(new_n634), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OR3_X1    g0710(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT109), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n910), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n673), .A2(G1), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n627), .A2(new_n900), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT44), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n627), .A2(new_n900), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT45), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n634), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n624), .B(new_n625), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n632), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n670), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n670), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n636), .B(KEYINPUT41), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n915), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n897), .B1(new_n914), .B2(new_n929), .ZN(G387));
  NOR2_X1   g0730(.A1(new_n394), .A2(G50), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT50), .ZN(new_n932));
  INV_X1    g0732(.A(new_n637), .ZN(new_n933));
  AOI211_X1 g0733(.A(G45), .B(new_n933), .C1(G68), .C2(G77), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n733), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n235), .B2(new_n734), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n738), .A2(new_n933), .B1(new_n437), .B2(new_n220), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n731), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n674), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT112), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n633), .A2(new_n896), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n701), .A2(G77), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n261), .C1(new_n440), .C2(new_n700), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n682), .B2(G150), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT113), .Z(new_n945));
  OAI22_X1  g0745(.A1(new_n202), .A2(new_n692), .B1(new_n689), .B2(new_n331), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n752), .A2(new_n277), .B1(new_n704), .B2(new_n392), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(G68), .C2(new_n696), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n261), .B1(new_n868), .B2(G116), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G317), .A2(new_n693), .B1(new_n690), .B2(G322), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n951), .B1(new_n697), .B2(new_n875), .C1(new_n754), .C2(new_n752), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT48), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n720), .A2(G283), .B1(G294), .B2(new_n701), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT49), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n950), .B1(new_n714), .B2(new_n681), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n949), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n940), .B(new_n941), .C1(new_n676), .C2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n925), .B2(new_n915), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n636), .B(KEYINPUT114), .Z(new_n964));
  NAND2_X1  g0764(.A1(new_n926), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n670), .A2(new_n925), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G393));
  NAND2_X1  g0767(.A1(new_n923), .A2(new_n926), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n964), .B1(new_n923), .B2(new_n926), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT116), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n923), .A2(new_n926), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT116), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n964), .A4(new_n968), .ZN(new_n974));
  INV_X1    g0774(.A(new_n915), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n923), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n903), .A2(new_n729), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n733), .A2(new_n246), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n730), .B1(new_n221), .B2(new_n440), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n675), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n704), .A2(new_n264), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n261), .B1(new_n508), .B2(new_n700), .C1(new_n697), .C2(new_n394), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(G50), .C2(new_n706), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n682), .A2(G143), .B1(G68), .B2(new_n701), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT115), .Z(new_n985));
  OAI22_X1  g0785(.A1(new_n763), .A2(new_n689), .B1(new_n692), .B2(new_n331), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT51), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G311), .A2(new_n693), .B1(new_n690), .B2(G317), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT52), .Z(new_n990));
  AOI21_X1  g0790(.A(new_n261), .B1(new_n868), .B2(G107), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n716), .B2(new_n702), .C1(new_n681), .C2(new_n717), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G116), .B2(new_n720), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G294), .A2(new_n696), .B1(new_n706), .B2(G303), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n980), .B1(new_n996), .B2(new_n676), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n976), .B1(new_n977), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n971), .A2(new_n974), .A3(new_n998), .ZN(G390));
  INV_X1    g0799(.A(KEYINPUT117), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n843), .ZN(new_n1001));
  OAI211_X1 g0801(.A(G330), .B(new_n773), .C1(new_n655), .C2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(new_n833), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(KEYINPUT117), .A3(new_n798), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n826), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n825), .B1(new_n807), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n824), .A2(new_n1007), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n616), .B1(new_n402), .B2(new_n771), .C1(new_n667), .C2(new_n668), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n769), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1009), .B1(new_n798), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1006), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1011), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1007), .B(new_n824), .C1(new_n1014), .C2(new_n833), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n660), .A2(new_n773), .A3(new_n798), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n826), .B1(new_n813), .B2(new_n798), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n825), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1013), .A2(new_n915), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(G128), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n689), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n701), .A2(G150), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT53), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(G125), .C2(new_n682), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT54), .B(G143), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT119), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n696), .A2(new_n1026), .B1(new_n706), .B2(G137), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n720), .A2(G159), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n261), .B1(new_n700), .B2(new_n202), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n693), .B2(G132), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n261), .B(new_n758), .C1(new_n682), .C2(G294), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n981), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n484), .A2(new_n692), .B1(new_n689), .B2(new_n716), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G87), .B2(new_n712), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G97), .A2(new_n696), .B1(new_n706), .B2(G107), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n749), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n674), .B(new_n1038), .C1(new_n277), .C2(new_n747), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n825), .B2(new_n728), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n405), .A2(G330), .A3(new_n849), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n838), .A2(new_n571), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n833), .B1(new_n659), .B2(new_n772), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1003), .A2(new_n1005), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n813), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1014), .B(new_n1016), .C1(new_n798), .C2(new_n1004), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1013), .A2(new_n1018), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(KEYINPUT118), .A3(new_n964), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1047), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT118), .B1(new_n1048), .B2(new_n964), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1019), .B(new_n1040), .C1(new_n1053), .C2(new_n1054), .ZN(G378));
  NAND3_X1  g0855(.A1(new_n846), .A2(new_n847), .A3(G330), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n291), .A2(new_n379), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n289), .A2(new_n613), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT122), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1056), .B(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n829), .B2(new_n836), .ZN(new_n1065));
  OAI21_X1  g0865(.A(KEYINPUT107), .B1(new_n816), .B2(new_n828), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n835), .A2(new_n830), .A3(new_n827), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n1063), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1042), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1065), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT57), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1065), .A2(KEYINPUT57), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n964), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n261), .A2(G41), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G50), .B(new_n1076), .C1(new_n257), .C2(new_n423), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n752), .A2(new_n440), .B1(new_n704), .B2(new_n312), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n700), .A2(new_n328), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n942), .A2(new_n1076), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n682), .C2(G283), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n437), .B2(new_n692), .C1(new_n484), .C2(new_n689), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1078), .B(new_n1082), .C1(new_n502), .C2(new_n696), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT120), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1077), .B1(new_n1084), .B2(KEYINPUT58), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1026), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1086), .A2(new_n702), .B1(new_n1020), .B2(new_n692), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n720), .A2(G150), .B1(G137), .B2(new_n696), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n760), .B2(new_n752), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(G125), .C2(new_n690), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n257), .B(new_n423), .C1(new_n700), .C2(new_n331), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n682), .B2(G124), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT59), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1085), .B1(KEYINPUT58), .B2(new_n1084), .C1(new_n1092), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n676), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT121), .Z(new_n1099));
  AOI211_X1 g0899(.A(new_n674), .B(new_n1099), .C1(new_n202), .C2(new_n747), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1061), .A2(new_n728), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1066), .A2(new_n1067), .A3(new_n1063), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1105), .B2(new_n915), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1075), .A2(new_n1106), .ZN(G375));
  NAND3_X1  g0907(.A1(new_n1045), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1051), .A2(new_n928), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n915), .B(KEYINPUT123), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n833), .A2(new_n727), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n676), .A2(G68), .A3(new_n727), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n712), .A2(G97), .B1(G283), .B2(new_n693), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n536), .B2(new_n689), .C1(new_n875), .C2(new_n681), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n720), .A2(new_n502), .B1(G116), .B2(new_n706), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n266), .B1(new_n700), .B2(new_n264), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT124), .Z(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(new_n437), .C2(new_n697), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n720), .A2(G50), .B1(G150), .B2(new_n696), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n266), .B(new_n1079), .C1(new_n690), .C2(G132), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n752), .C2(new_n1086), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n682), .A2(G128), .B1(G137), .B2(new_n693), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n712), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n331), .B2(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1115), .A2(new_n1119), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n674), .B(new_n1113), .C1(new_n1126), .C2(new_n676), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1110), .A2(new_n1111), .B1(new_n1112), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1109), .A2(new_n1128), .ZN(G381));
  INV_X1    g0929(.A(G378), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1075), .A2(new_n1130), .A3(new_n1106), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(G387), .A2(G390), .ZN(new_n1133));
  NOR4_X1   g0933(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(G407));
  OAI211_X1 g0935(.A(G407), .B(G213), .C1(G343), .C2(new_n1131), .ZN(G409));
  AOI21_X1  g0936(.A(KEYINPUT57), .B1(new_n1105), .B2(new_n1070), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1074), .A2(new_n964), .ZN(new_n1138));
  OAI211_X1 g0938(.A(G378), .B(new_n1106), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1102), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1111), .B1(new_n1070), .B2(new_n928), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1130), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n614), .A2(G213), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n964), .B(new_n1051), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1128), .ZN(new_n1150));
  INV_X1    g0950(.A(G384), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(G384), .A3(new_n1128), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1145), .A2(new_n1146), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT62), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1146), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(G2897), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(G2897), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1152), .A2(new_n1153), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT61), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT62), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1145), .A2(new_n1166), .A3(new_n1146), .A4(new_n1155), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1157), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1133), .ZN(new_n1169));
  XOR2_X1   g0969(.A(G393), .B(G396), .Z(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(G387), .A2(G390), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(G387), .A2(G390), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1170), .B1(new_n1174), .B2(new_n1133), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1168), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT63), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1156), .B1(new_n1163), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1173), .A2(new_n1175), .A3(new_n1165), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1158), .B(new_n1154), .C1(new_n1139), .C2(new_n1144), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(KEYINPUT63), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1179), .A2(new_n1182), .A3(KEYINPUT125), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT125), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(G405));
  INV_X1    g0985(.A(new_n1176), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1139), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G378), .B1(new_n1075), .B2(new_n1106), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT126), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1154), .A2(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1154), .A2(KEYINPUT127), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1188), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(KEYINPUT126), .A3(new_n1139), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(new_n1176), .A3(new_n1192), .A4(new_n1191), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(G402));
endmodule


