//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT79), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G155gat), .B(G162gat), .ZN(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  INV_X1    g019(.A(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT2), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  AND2_X1   g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT22), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n231));
  INV_X1    g030(.A(G204gat), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n234));
  AOI21_X1  g033(.A(G204gat), .B1(new_n234), .B2(new_n229), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n228), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI221_X1 g038(.A(new_n228), .B1(new_n226), .B2(new_n237), .C1(new_n233), .C2(new_n235), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT29), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT81), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n225), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI211_X1 g042(.A(KEYINPUT81), .B(KEYINPUT29), .C1(new_n239), .C2(new_n240), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n224), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n240), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n223), .A3(new_n225), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n213), .A2(new_n223), .A3(KEYINPUT76), .A4(new_n225), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G228gat), .A2(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n224), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n232), .B1(new_n230), .B2(new_n231), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n234), .A2(G204gat), .A3(new_n229), .ZN(new_n259));
  AOI211_X1 g058(.A(new_n227), .B(new_n238), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT29), .B1(new_n260), .B2(KEYINPUT80), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n239), .A2(new_n240), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n257), .B1(new_n264), .B2(new_n225), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n254), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n206), .B1(new_n256), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n256), .A2(new_n266), .A3(new_n206), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI211_X1 g069(.A(KEYINPUT82), .B(new_n206), .C1(new_n256), .C2(new_n266), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n205), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n267), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n269), .A3(new_n204), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276));
  INV_X1    g075(.A(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G113gat), .ZN(new_n278));
  INV_X1    g077(.A(G113gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G120gat), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT1), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G127gat), .B(G134gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(G127gat), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(G134gat), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n281), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n287), .A2(new_n292), .A3(KEYINPUT72), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n276), .B1(new_n297), .B2(new_n224), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n287), .A2(new_n292), .A3(KEYINPUT72), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT72), .B1(new_n287), .B2(new_n292), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n299), .A2(new_n300), .A3(new_n281), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT4), .B(new_n257), .C1(new_n301), .C2(new_n284), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n308), .B2(new_n251), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT5), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n285), .A2(G127gat), .A3(new_n286), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n315));
  INV_X1    g114(.A(G134gat), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n294), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n281), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n296), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n320), .A2(new_n224), .A3(new_n283), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n224), .B1(new_n320), .B2(new_n283), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n306), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n304), .A2(new_n309), .B1(KEYINPUT77), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n257), .B1(new_n301), .B2(new_n284), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n224), .A3(new_n283), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n305), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT78), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n251), .A2(new_n297), .A3(new_n307), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n305), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n303), .A2(new_n333), .B1(new_n328), .B2(new_n329), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT5), .B1(new_n323), .B2(KEYINPUT77), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n312), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT6), .ZN(new_n343));
  INV_X1    g142(.A(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT6), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n336), .B1(new_n334), .B2(new_n335), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n310), .A2(new_n330), .A3(KEYINPUT78), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n311), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n345), .A3(new_n344), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n275), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n246), .ZN(new_n356));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G169gat), .ZN(new_n359));
  INV_X1    g158(.A(G176gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT23), .ZN(new_n361));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT64), .B1(new_n364), .B2(KEYINPUT23), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(new_n360), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT66), .B(G190gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT65), .B(G183gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT24), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(G183gat), .A3(G190gat), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n371), .A2(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n377), .B2(KEYINPUT67), .ZN(new_n378));
  INV_X1    g177(.A(G190gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT66), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT66), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(G183gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT65), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G183gat), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n380), .A2(new_n382), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n374), .A2(new_n376), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n387), .A2(KEYINPUT67), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT25), .B1(new_n378), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n364), .A2(new_n391), .B1(new_n362), .B2(KEYINPUT69), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n393));
  NOR4_X1   g192(.A1(new_n393), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT68), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n395), .A2(new_n397), .B1(G183gat), .B2(G190gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n372), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT28), .B1(new_n402), .B2(new_n371), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT27), .B(G183gat), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n371), .A2(new_n404), .A3(KEYINPUT28), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n370), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n358), .B1(new_n410), .B2(new_n252), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n370), .A2(new_n407), .A3(new_n408), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n401), .B1(new_n384), .B2(new_n386), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n371), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT28), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n405), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n412), .B1(new_n418), .B2(new_n398), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n357), .B1(new_n419), .B2(new_n390), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n356), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n422));
  NOR3_X1   g221(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT69), .ZN(new_n424));
  AND2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n393), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n424), .B1(new_n426), .B2(new_n423), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n396), .B(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n373), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n409), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT67), .B1(new_n387), .B2(new_n388), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n425), .B1(KEYINPUT23), .B2(new_n364), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n364), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n377), .A2(KEYINPUT67), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n407), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n252), .B1(new_n431), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n357), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n410), .A2(new_n358), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n246), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND3_X1  g245(.A1(new_n421), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT30), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n446), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n411), .A2(new_n356), .A3(new_n420), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n246), .B1(new_n441), .B2(new_n442), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n297), .B1(new_n431), .B2(new_n439), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n320), .A2(new_n283), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n390), .A2(new_n406), .A3(new_n459), .A4(new_n409), .ZN(new_n460));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT34), .Z(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n458), .B2(new_n460), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT33), .ZN(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G43gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G71gat), .B(G99gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n458), .A2(new_n460), .ZN(new_n471));
  INV_X1    g270(.A(new_n461), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n468), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT73), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n479));
  NOR4_X1   g278(.A1(new_n464), .A2(new_n479), .A3(new_n469), .A4(new_n476), .ZN(new_n480));
  OAI221_X1 g279(.A(new_n463), .B1(new_n465), .B2(new_n470), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n478), .A2(new_n480), .B1(new_n465), .B2(new_n470), .ZN(new_n482));
  INV_X1    g281(.A(new_n463), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n457), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n355), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n482), .B2(KEYINPUT74), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n483), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n275), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n353), .A2(new_n457), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT35), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n482), .A2(KEYINPUT74), .A3(new_n483), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT36), .B1(new_n494), .B2(new_n487), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n484), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n338), .A2(new_n344), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n332), .A2(new_n298), .A3(new_n302), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT39), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n306), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n342), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n326), .A2(new_n305), .A3(new_n327), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT39), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n306), .B2(new_n500), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT84), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT40), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n500), .A2(new_n306), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n321), .A2(new_n322), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n510), .B2(new_n305), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n342), .A3(new_n502), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT84), .B1(new_n513), .B2(KEYINPUT83), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT84), .B(KEYINPUT40), .C1(new_n513), .C2(KEYINPUT83), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n456), .B(new_n499), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT38), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n453), .B2(new_n454), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n421), .A2(new_n443), .A3(KEYINPUT38), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n448), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n519), .B(new_n520), .C1(KEYINPUT37), .C2(new_n446), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n347), .A2(new_n523), .A3(new_n352), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(new_n525), .A3(new_n275), .ZN(new_n526));
  INV_X1    g325(.A(new_n275), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n491), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n498), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n493), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT95), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534));
  AND2_X1   g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT9), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n532), .A2(new_n536), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n534), .A2(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(KEYINPUT94), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n546), .B(new_n547), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(new_n289), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(G1gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT16), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(G1gat), .B2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G8gat), .ZN(new_n555));
  INV_X1    g354(.A(G8gat), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n553), .B(new_n556), .C1(G1gat), .C2(new_n550), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n545), .B2(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n548), .B(G127gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n559), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(new_n220), .ZN(new_n565));
  XOR2_X1   g364(.A(G183gat), .B(G211gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n560), .B2(new_n563), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n573), .A2(KEYINPUT8), .ZN(new_n574));
  NOR2_X1   g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(KEYINPUT8), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(KEYINPUT97), .C1(G85gat), .C2(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(G85gat), .A3(G92gat), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n580), .A3(new_n581), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G99gat), .B(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT98), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n586), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n578), .B2(new_n576), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT99), .B1(new_n593), .B2(new_n589), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n588), .A2(new_n598), .A3(new_n590), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(G29gat), .A2(G36gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT14), .ZN(new_n602));
  XOR2_X1   g401(.A(G43gat), .B(G50gat), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT15), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT89), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT88), .B(G36gat), .Z(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(G29gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n609), .A3(G29gat), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n606), .A2(new_n608), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n602), .A3(new_n605), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n607), .B1(new_n615), .B2(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n616), .A3(KEYINPUT17), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n600), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n600), .ZN(new_n624));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625));
  AND2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n626), .B2(new_n627), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n571), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n637));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n618), .B2(new_n558), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n641), .A3(new_n558), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n618), .A2(new_n558), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n555), .A2(new_n557), .A3(KEYINPUT90), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT90), .B1(new_n555), .B2(new_n557), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n620), .A2(new_n617), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n644), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n651), .B(new_n638), .C1(new_n652), .C2(new_n642), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT92), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n647), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT18), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n653), .A2(KEYINPUT92), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G113gat), .B(G141gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G169gat), .B(G197gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n655), .A2(new_n667), .A3(new_n657), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n588), .A2(KEYINPUT98), .A3(new_n590), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n594), .B1(new_n593), .B2(new_n589), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n597), .A2(new_n599), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n544), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT10), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n588), .A2(KEYINPUT100), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n588), .A2(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n590), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n596), .B(new_n545), .C1(new_n679), .C2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n677), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n544), .A2(new_n678), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n596), .A2(new_n597), .A3(new_n599), .A4(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n672), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n671), .B1(new_n677), .B2(new_n682), .ZN(new_n687));
  XOR2_X1   g486(.A(G120gat), .B(G148gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT101), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n686), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n686), .B2(new_n687), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n636), .A2(new_n670), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n530), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n353), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(new_n551), .ZN(G1324gat));
  INV_X1    g498(.A(new_n697), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n556), .B1(new_n700), .B2(new_n456), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT16), .B(G8gat), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n697), .A2(new_n457), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT42), .B2(new_n703), .ZN(G1325gat));
  OAI21_X1  g504(.A(G15gat), .B1(new_n697), .B2(new_n498), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n481), .A2(new_n484), .ZN(new_n707));
  INV_X1    g506(.A(G15gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n697), .B2(new_n709), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n697), .A2(new_n275), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(G29gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n353), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n571), .A2(new_n670), .A3(new_n695), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT102), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n634), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n456), .B1(new_n347), .B2(new_n352), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n495), .B(new_n497), .C1(new_n275), .C2(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n517), .A2(new_n525), .A3(new_n275), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT103), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n498), .A2(new_n724), .A3(new_n526), .A4(new_n528), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n719), .B1(new_n726), .B2(new_n493), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n718), .B1(new_n530), .B2(new_n634), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n715), .B(new_n717), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n714), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n530), .A2(new_n634), .A3(new_n716), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n714), .A3(new_n715), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(G1328gat));
  OR2_X1    g536(.A1(new_n727), .A2(new_n728), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n456), .A3(new_n717), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n610), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n733), .A2(new_n457), .A3(new_n610), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1329gat));
  INV_X1    g542(.A(G43gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n498), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(new_n717), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n734), .A2(new_n707), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n747), .A2(new_n744), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n748));
  OR2_X1    g547(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n746), .B2(new_n748), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(G1330gat));
  AND2_X1   g551(.A1(new_n527), .A2(G50gat), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n738), .A2(new_n717), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n275), .B1(new_n733), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(G50gat), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT48), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n758), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n738), .A2(new_n717), .A3(new_n753), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(G1331gat));
  NAND4_X1  g563(.A1(new_n720), .A2(new_n275), .A3(new_n488), .A4(new_n489), .ZN(new_n765));
  AOI22_X1  g564(.A1(KEYINPUT35), .A2(new_n765), .B1(new_n355), .B2(new_n485), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n723), .B2(new_n725), .ZN(new_n767));
  INV_X1    g566(.A(new_n695), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n767), .A2(new_n669), .A3(new_n636), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n715), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT107), .B(G57gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n456), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT49), .B(G64gat), .Z(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(G1333gat));
  INV_X1    g575(.A(new_n498), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n769), .A2(G71gat), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n707), .B(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(G71gat), .B1(new_n769), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT50), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n769), .A2(new_n782), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(new_n778), .C1(new_n786), .C2(G71gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n527), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g589(.A1(new_n571), .A2(new_n669), .A3(new_n768), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n738), .A2(new_n715), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G85gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n570), .A2(new_n670), .A3(new_n634), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n726), .B2(new_n493), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n726), .A2(new_n493), .ZN(new_n797));
  INV_X1    g596(.A(new_n794), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT51), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n795), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OR3_X1    g602(.A1(new_n353), .A2(new_n768), .A3(G85gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n793), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  OAI211_X1 g604(.A(new_n456), .B(new_n791), .C1(new_n727), .C2(new_n728), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n806), .B2(G92gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n768), .A2(new_n457), .A3(G92gat), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n767), .B2(new_n794), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT109), .B1(new_n795), .B2(KEYINPUT51), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n767), .A2(new_n800), .A3(new_n814), .A4(new_n794), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n816), .A2(new_n808), .B1(G92gat), .B2(new_n806), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n810), .B1(new_n817), .B2(new_n818), .ZN(G1337gat));
  INV_X1    g618(.A(G99gat), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n777), .B(new_n791), .C1(new_n727), .C2(new_n728), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n707), .A2(new_n820), .A3(new_n695), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n825), .B(KEYINPUT112), .Z(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n803), .B2(new_n826), .ZN(G1338gat));
  XNOR2_X1  g626(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n527), .B(new_n791), .C1(new_n727), .C2(new_n728), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(G106gat), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n275), .A2(new_n768), .A3(G106gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n803), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n831), .B(KEYINPUT113), .Z(new_n833));
  AOI22_X1  g632(.A1(new_n816), .A2(new_n833), .B1(G106gat), .B2(new_n829), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n683), .A2(new_n685), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n671), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n692), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n685), .A2(new_n672), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n683), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n686), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n837), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n686), .A2(new_n687), .A3(new_n692), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n671), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n683), .B2(new_n842), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n837), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n691), .B1(new_n686), .B2(new_n839), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n657), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n656), .B1(new_n653), .B2(KEYINPUT92), .ZN(new_n855));
  NOR4_X1   g654(.A1(new_n854), .A2(new_n855), .A3(new_n665), .A4(new_n647), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n667), .B1(new_n655), .B2(new_n657), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n846), .B(new_n853), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n663), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n645), .A2(new_n651), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(G229gat), .A3(G233gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n645), .A2(new_n646), .A3(new_n640), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n859), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n695), .A3(new_n668), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n634), .B1(new_n858), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n867), .A2(new_n632), .A3(new_n668), .A4(new_n633), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n853), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n570), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n571), .A2(new_n670), .A3(new_n635), .A4(new_n768), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n353), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n456), .A3(new_n490), .ZN(new_n877));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n669), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n874), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n485), .A2(new_n275), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n715), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n875), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n670), .A2(new_n279), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(G1340gat));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n695), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G120gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n877), .A2(new_n277), .A3(new_n695), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1341gat));
  NAND2_X1  g694(.A1(new_n885), .A2(new_n571), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n315), .B2(new_n314), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n290), .A3(new_n291), .A4(new_n571), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1342gat));
  NOR2_X1   g698(.A1(new_n876), .A2(new_n490), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n635), .A2(new_n456), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n285), .A3(new_n286), .A4(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n885), .A2(new_n634), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n316), .ZN(G1343gat));
  NAND3_X1  g705(.A1(new_n498), .A2(new_n715), .A3(new_n457), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n275), .B1(new_n873), .B2(new_n874), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT55), .B1(new_n844), .B2(new_n686), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n693), .B1(new_n912), .B2(new_n841), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n848), .A2(new_n850), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT55), .B1(new_n914), .B2(new_n852), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n846), .A2(new_n853), .A3(KEYINPUT119), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n669), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n634), .B1(new_n918), .B2(new_n868), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n570), .B1(new_n919), .B2(new_n872), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n275), .B1(new_n920), .B2(new_n874), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n910), .B(new_n669), .C1(new_n921), .C2(new_n909), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G141gat), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n498), .A2(new_n527), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n925), .A2(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(KEYINPUT121), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n875), .A2(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n670), .A2(G141gat), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n457), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n923), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT58), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1344gat));
  AND3_X1   g735(.A1(new_n928), .A2(new_n929), .A3(new_n457), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n216), .A3(new_n695), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n910), .B1(new_n921), .B2(new_n909), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n768), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G148gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n909), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n908), .A2(new_n909), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n907), .A2(new_n768), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n938), .B1(new_n943), .B2(new_n948), .ZN(G1345gat));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n220), .A3(new_n571), .ZN(new_n950));
  OAI21_X1  g749(.A(G155gat), .B1(new_n939), .B2(new_n570), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1346gat));
  OAI21_X1  g751(.A(G162gat), .B1(new_n939), .B2(new_n635), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n928), .A2(new_n929), .A3(new_n221), .A4(new_n901), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1347gat));
  NAND2_X1  g754(.A1(new_n353), .A2(new_n456), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n781), .A2(new_n527), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n879), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n879), .A2(new_n957), .A3(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n359), .A3(new_n670), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n715), .B1(new_n873), .B2(new_n874), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n490), .A2(new_n457), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n669), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n963), .A2(new_n968), .ZN(G1348gat));
  NOR3_X1   g768(.A1(new_n962), .A2(new_n360), .A3(new_n768), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n360), .B1(new_n966), .B2(new_n768), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(G1349gat));
  INV_X1    g774(.A(new_n372), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n976), .B1(new_n962), .B2(new_n570), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n967), .A2(new_n404), .A3(new_n571), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT60), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n960), .A2(new_n634), .A3(new_n961), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G190gat), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(KEYINPUT61), .A3(new_n988), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n967), .A2(new_n371), .A3(new_n634), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT124), .B1(new_n984), .B2(G190gat), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n989), .A2(new_n993), .ZN(G1351gat));
  AND2_X1   g793(.A1(new_n944), .A2(new_n945), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n777), .A2(new_n956), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n996), .B(KEYINPUT126), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(G197gat), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n670), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n925), .A2(new_n457), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n964), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n964), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1004), .A2(new_n669), .A3(new_n1006), .ZN(new_n1007));
  AOI22_X1  g806(.A1(new_n999), .A2(new_n1001), .B1(new_n1000), .B2(new_n1007), .ZN(G1352gat));
  OAI21_X1  g807(.A(G204gat), .B1(new_n998), .B2(new_n768), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1003), .A2(G204gat), .A3(new_n768), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1353gat));
  NAND4_X1  g811(.A1(new_n944), .A2(new_n571), .A3(new_n945), .A4(new_n997), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(G211gat), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(KEYINPUT63), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT63), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1013), .A2(new_n1016), .A3(G211gat), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n570), .A2(G211gat), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1004), .A2(new_n1006), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(KEYINPUT127), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1021));
  NAND4_X1  g820(.A1(new_n1004), .A2(new_n1021), .A3(new_n1006), .A4(new_n1018), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1015), .A2(new_n1017), .A3(new_n1023), .ZN(G1354gat));
  OAI21_X1  g823(.A(G218gat), .B1(new_n998), .B2(new_n635), .ZN(new_n1025));
  NOR2_X1   g824(.A1(new_n635), .A2(G218gat), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1004), .A2(new_n1006), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1025), .A2(new_n1027), .ZN(G1355gat));
endmodule


