

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n770), .B(KEYINPUT32), .ZN(n799) );
  NOR2_X4 U552 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  NOR2_X1 U553 ( .A1(n717), .A2(n950), .ZN(n719) );
  NOR2_X1 U554 ( .A1(n755), .A2(n712), .ZN(n714) );
  BUF_X1 U555 ( .A(n613), .Z(n614) );
  INV_X1 U556 ( .A(KEYINPUT64), .ZN(n789) );
  NOR2_X1 U557 ( .A1(G651), .A2(n651), .ZN(n646) );
  NOR2_X2 U558 ( .A1(n651), .A2(n536), .ZN(n555) );
  NOR2_X1 U559 ( .A1(n795), .A2(n794), .ZN(n515) );
  INV_X1 U560 ( .A(KEYINPUT66), .ZN(n718) );
  XNOR2_X1 U561 ( .A(n719), .B(n718), .ZN(n727) );
  XNOR2_X1 U562 ( .A(n762), .B(KEYINPUT102), .ZN(n763) );
  XNOR2_X1 U563 ( .A(n764), .B(n763), .ZN(n773) );
  AND2_X1 U564 ( .A1(n769), .A2(n768), .ZN(n770) );
  INV_X1 U565 ( .A(n961), .ZN(n794) );
  NAND2_X1 U566 ( .A1(n711), .A2(n710), .ZN(n755) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n679) );
  XOR2_X1 U568 ( .A(KEYINPUT65), .B(n679), .Z(n711) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n517) );
  NOR2_X2 U570 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U571 ( .A1(n867), .A2(G137), .ZN(n528) );
  NOR2_X1 U572 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U573 ( .A(KEYINPUT76), .B(n562), .Z(n950) );
  NOR2_X1 U574 ( .A1(n533), .A2(n532), .ZN(G160) );
  INV_X1 U575 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n521), .A2(G2104), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n516), .B(KEYINPUT67), .ZN(n613) );
  NAND2_X1 U578 ( .A1(G102), .A2(n613), .ZN(n520) );
  XNOR2_X2 U579 ( .A(n518), .B(n517), .ZN(n867) );
  NAND2_X1 U580 ( .A1(G138), .A2(n867), .ZN(n519) );
  NAND2_X1 U581 ( .A1(n520), .A2(n519), .ZN(n525) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U583 ( .A1(G114), .A2(n870), .ZN(n523) );
  NOR2_X2 U584 ( .A1(G2104), .A2(n521), .ZN(n872) );
  NAND2_X1 U585 ( .A1(G126), .A2(n872), .ZN(n522) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n525), .A2(n524), .ZN(G164) );
  NAND2_X1 U588 ( .A1(G113), .A2(n870), .ZN(n527) );
  NAND2_X1 U589 ( .A1(G125), .A2(n872), .ZN(n526) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n533) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT68), .ZN(n531) );
  NAND2_X1 U592 ( .A1(G101), .A2(n613), .ZN(n529) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U595 ( .A(G651), .ZN(n536) );
  NOR2_X1 U596 ( .A1(G543), .A2(n536), .ZN(n534) );
  XOR2_X2 U597 ( .A(KEYINPUT1), .B(n534), .Z(n650) );
  NAND2_X1 U598 ( .A1(G64), .A2(n650), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT69), .ZN(n542) );
  XOR2_X1 U600 ( .A(G543), .B(KEYINPUT0), .Z(n651) );
  NAND2_X1 U601 ( .A1(n555), .A2(G77), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT70), .ZN(n539) );
  NAND2_X1 U603 ( .A1(G90), .A2(n638), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n646), .A2(G52), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(G301) );
  INV_X1 U609 ( .A(G301), .ZN(G171) );
  NAND2_X1 U610 ( .A1(G60), .A2(n650), .ZN(n546) );
  NAND2_X1 U611 ( .A1(G47), .A2(n646), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U613 ( .A1(G85), .A2(n638), .ZN(n548) );
  NAND2_X1 U614 ( .A1(G72), .A2(n555), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(G290) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G860), .ZN(n606) );
  NAND2_X1 U619 ( .A1(n650), .A2(G56), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n551), .B(KEYINPUT14), .ZN(n553) );
  NAND2_X1 U621 ( .A1(G43), .A2(n646), .ZN(n552) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n638), .A2(G81), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n554), .B(KEYINPUT12), .ZN(n557) );
  NAND2_X1 U625 ( .A1(G68), .A2(n555), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(KEYINPUT75), .B(n558), .ZN(n559) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(n559), .ZN(n560) );
  OR2_X1 U629 ( .A1(n606), .A2(n950), .ZN(G153) );
  NAND2_X1 U630 ( .A1(n646), .A2(G50), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G88), .A2(n638), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G75), .A2(n555), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n650), .A2(G62), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT88), .B(n565), .Z(n566) );
  NOR2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT89), .B(n570), .Z(G303) );
  INV_X1 U639 ( .A(G303), .ZN(G166) );
  INV_X1 U640 ( .A(G132), .ZN(G219) );
  INV_X1 U641 ( .A(G82), .ZN(G220) );
  NAND2_X1 U642 ( .A1(n555), .A2(G76), .ZN(n571) );
  XNOR2_X1 U643 ( .A(KEYINPUT78), .B(n571), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n638), .A2(G89), .ZN(n572) );
  XNOR2_X1 U645 ( .A(KEYINPUT4), .B(n572), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U647 ( .A(n575), .B(KEYINPUT5), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G63), .A2(n650), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G51), .A2(n646), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U651 ( .A(KEYINPUT6), .B(n578), .Z(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U654 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n582), .B(KEYINPUT10), .ZN(n583) );
  XNOR2_X1 U657 ( .A(KEYINPUT74), .B(n583), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n830) );
  NAND2_X1 U659 ( .A1(n830), .A2(G567), .ZN(n584) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G92), .A2(n638), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G66), .A2(n650), .ZN(n586) );
  NAND2_X1 U664 ( .A1(G54), .A2(n646), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U666 ( .A1(G79), .A2(n555), .ZN(n587) );
  XNOR2_X1 U667 ( .A(KEYINPUT77), .B(n587), .ZN(n588) );
  NOR2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT15), .ZN(n943) );
  INV_X1 U671 ( .A(n943), .ZN(n726) );
  INV_X1 U672 ( .A(G868), .ZN(n663) );
  NAND2_X1 U673 ( .A1(n726), .A2(n663), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G53), .A2(n646), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n595), .B(KEYINPUT72), .ZN(n602) );
  NAND2_X1 U677 ( .A1(G91), .A2(n638), .ZN(n597) );
  NAND2_X1 U678 ( .A1(G78), .A2(n555), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U680 ( .A1(G65), .A2(n650), .ZN(n598) );
  XNOR2_X1 U681 ( .A(KEYINPUT71), .B(n598), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(G299) );
  NOR2_X1 U684 ( .A1(G286), .A2(n663), .ZN(n603) );
  XOR2_X1 U685 ( .A(KEYINPUT79), .B(n603), .Z(n605) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n607), .A2(n943), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n608), .B(KEYINPUT80), .ZN(n609) );
  XNOR2_X1 U691 ( .A(KEYINPUT16), .B(n609), .ZN(G148) );
  NOR2_X1 U692 ( .A1(n950), .A2(G868), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G868), .A2(n943), .ZN(n610) );
  NOR2_X1 U694 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U695 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G99), .A2(n614), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G111), .A2(n870), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n872), .A2(G123), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT18), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G135), .A2(n867), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U703 ( .A(KEYINPUT81), .B(n620), .Z(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n1001) );
  XOR2_X1 U705 ( .A(G2096), .B(n1001), .Z(n623) );
  NOR2_X1 U706 ( .A1(G2100), .A2(n623), .ZN(n624) );
  XOR2_X1 U707 ( .A(KEYINPUT82), .B(n624), .Z(G156) );
  NAND2_X1 U708 ( .A1(G80), .A2(n555), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n625), .B(KEYINPUT84), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G67), .A2(n650), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G55), .A2(n646), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G93), .A2(n638), .ZN(n628) );
  XNOR2_X1 U714 ( .A(KEYINPUT83), .B(n628), .ZN(n629) );
  NOR2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n664) );
  NAND2_X1 U717 ( .A1(G559), .A2(n943), .ZN(n633) );
  XNOR2_X1 U718 ( .A(n633), .B(n950), .ZN(n660) );
  NOR2_X1 U719 ( .A1(G860), .A2(n660), .ZN(n634) );
  XNOR2_X1 U720 ( .A(n634), .B(KEYINPUT85), .ZN(n635) );
  XNOR2_X1 U721 ( .A(n664), .B(n635), .ZN(G145) );
  XOR2_X1 U722 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n637) );
  NAND2_X1 U723 ( .A1(G73), .A2(n555), .ZN(n636) );
  XNOR2_X1 U724 ( .A(n637), .B(n636), .ZN(n642) );
  NAND2_X1 U725 ( .A1(G61), .A2(n650), .ZN(n640) );
  NAND2_X1 U726 ( .A1(G86), .A2(n638), .ZN(n639) );
  NAND2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U729 ( .A(KEYINPUT87), .B(n643), .Z(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(G48), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G49), .A2(n646), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U736 ( .A1(n651), .A2(G87), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n653), .A2(n652), .ZN(G288) );
  XOR2_X1 U738 ( .A(G290), .B(G305), .Z(n654) );
  XNOR2_X1 U739 ( .A(n664), .B(n654), .ZN(n657) );
  XOR2_X1 U740 ( .A(KEYINPUT90), .B(KEYINPUT19), .Z(n655) );
  XNOR2_X1 U741 ( .A(G288), .B(n655), .ZN(n656) );
  XOR2_X1 U742 ( .A(n657), .B(n656), .Z(n659) );
  INV_X1 U743 ( .A(G299), .ZN(n738) );
  XNOR2_X1 U744 ( .A(n738), .B(G166), .ZN(n658) );
  XNOR2_X1 U745 ( .A(n659), .B(n658), .ZN(n886) );
  XNOR2_X1 U746 ( .A(n886), .B(n660), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n661), .A2(G868), .ZN(n662) );
  XOR2_X1 U748 ( .A(KEYINPUT91), .B(n662), .Z(n666) );
  NAND2_X1 U749 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n667) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U758 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U759 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G69), .A2(n672), .ZN(n917) );
  NAND2_X1 U761 ( .A1(n917), .A2(G567), .ZN(n677) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U764 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U765 ( .A1(G96), .A2(n675), .ZN(n918) );
  NAND2_X1 U766 ( .A1(n918), .A2(G2106), .ZN(n676) );
  NAND2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n844) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U769 ( .A1(n844), .A2(n678), .ZN(n833) );
  NAND2_X1 U770 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n709) );
  NOR2_X1 U772 ( .A1(n711), .A2(n709), .ZN(n825) );
  XOR2_X1 U773 ( .A(G2067), .B(KEYINPUT37), .Z(n680) );
  XOR2_X1 U774 ( .A(KEYINPUT92), .B(n680), .Z(n823) );
  NAND2_X1 U775 ( .A1(G104), .A2(n614), .ZN(n682) );
  NAND2_X1 U776 ( .A1(G140), .A2(n867), .ZN(n681) );
  NAND2_X1 U777 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U778 ( .A(KEYINPUT34), .B(n683), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G116), .A2(n870), .ZN(n685) );
  NAND2_X1 U780 ( .A1(G128), .A2(n872), .ZN(n684) );
  NAND2_X1 U781 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U782 ( .A(n686), .B(KEYINPUT35), .Z(n687) );
  NOR2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U784 ( .A(KEYINPUT36), .B(n689), .Z(n690) );
  XNOR2_X1 U785 ( .A(KEYINPUT93), .B(n690), .ZN(n883) );
  OR2_X1 U786 ( .A1(n823), .A2(n883), .ZN(n691) );
  XNOR2_X1 U787 ( .A(n691), .B(KEYINPUT94), .ZN(n821) );
  NAND2_X1 U788 ( .A1(G95), .A2(n614), .ZN(n693) );
  NAND2_X1 U789 ( .A1(G107), .A2(n870), .ZN(n692) );
  NAND2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U791 ( .A1(G131), .A2(n867), .ZN(n695) );
  NAND2_X1 U792 ( .A1(G119), .A2(n872), .ZN(n694) );
  NAND2_X1 U793 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n852) );
  NAND2_X1 U795 ( .A1(G1991), .A2(n852), .ZN(n698) );
  XNOR2_X1 U796 ( .A(n698), .B(KEYINPUT95), .ZN(n707) );
  NAND2_X1 U797 ( .A1(G117), .A2(n870), .ZN(n700) );
  NAND2_X1 U798 ( .A1(G129), .A2(n872), .ZN(n699) );
  NAND2_X1 U799 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n614), .A2(G105), .ZN(n701) );
  XOR2_X1 U801 ( .A(KEYINPUT38), .B(n701), .Z(n702) );
  NOR2_X1 U802 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n867), .A2(G141), .ZN(n704) );
  NAND2_X1 U804 ( .A1(n705), .A2(n704), .ZN(n880) );
  AND2_X1 U805 ( .A1(G1996), .A2(n880), .ZN(n706) );
  NOR2_X1 U806 ( .A1(n707), .A2(n706), .ZN(n816) );
  NAND2_X1 U807 ( .A1(n821), .A2(n816), .ZN(n1015) );
  NAND2_X1 U808 ( .A1(n825), .A2(n1015), .ZN(n708) );
  XOR2_X1 U809 ( .A(KEYINPUT96), .B(n708), .Z(n812) );
  INV_X1 U810 ( .A(n709), .ZN(n710) );
  INV_X1 U811 ( .A(G1996), .ZN(n712) );
  XNOR2_X1 U812 ( .A(KEYINPUT26), .B(KEYINPUT99), .ZN(n713) );
  XNOR2_X1 U813 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n755), .A2(G1341), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n716), .A2(n715), .ZN(n717) );
  INV_X1 U816 ( .A(n727), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n720), .A2(n943), .ZN(n724) );
  INV_X1 U818 ( .A(n755), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n744), .A2(G1348), .ZN(n722) );
  NOR2_X1 U820 ( .A1(G2067), .A2(n755), .ZN(n721) );
  NOR2_X1 U821 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U823 ( .A(n725), .B(KEYINPUT100), .ZN(n729) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n736) );
  INV_X1 U826 ( .A(G2072), .ZN(n996) );
  NOR2_X1 U827 ( .A1(n755), .A2(n996), .ZN(n731) );
  XOR2_X1 U828 ( .A(KEYINPUT27), .B(KEYINPUT97), .Z(n730) );
  XNOR2_X1 U829 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U830 ( .A1(n755), .A2(G1956), .ZN(n732) );
  NAND2_X1 U831 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U832 ( .A(KEYINPUT98), .B(n734), .Z(n737) );
  NAND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n735) );
  NAND2_X1 U834 ( .A1(n736), .A2(n735), .ZN(n741) );
  NOR2_X1 U835 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U836 ( .A(n739), .B(KEYINPUT28), .Z(n740) );
  NAND2_X1 U837 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U838 ( .A(KEYINPUT101), .B(KEYINPUT29), .ZN(n742) );
  XNOR2_X1 U839 ( .A(n743), .B(n742), .ZN(n771) );
  INV_X1 U840 ( .A(G1961), .ZN(n919) );
  NAND2_X1 U841 ( .A1(n755), .A2(n919), .ZN(n746) );
  XNOR2_X1 U842 ( .A(KEYINPUT25), .B(G2078), .ZN(n970) );
  NAND2_X1 U843 ( .A1(n744), .A2(n970), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n746), .A2(n745), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n759), .A2(G171), .ZN(n772) );
  NAND2_X1 U846 ( .A1(G8), .A2(n755), .ZN(n806) );
  NOR2_X1 U847 ( .A1(G1971), .A2(n806), .ZN(n748) );
  NOR2_X1 U848 ( .A1(G2090), .A2(n755), .ZN(n747) );
  NOR2_X1 U849 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U850 ( .A(KEYINPUT103), .B(n749), .Z(n750) );
  NAND2_X1 U851 ( .A1(n750), .A2(G303), .ZN(n765) );
  INV_X1 U852 ( .A(n765), .ZN(n751) );
  OR2_X1 U853 ( .A1(n751), .A2(G286), .ZN(n752) );
  AND2_X1 U854 ( .A1(G8), .A2(n752), .ZN(n754) );
  AND2_X1 U855 ( .A1(n772), .A2(n754), .ZN(n753) );
  NAND2_X1 U856 ( .A1(n771), .A2(n753), .ZN(n769) );
  INV_X1 U857 ( .A(n754), .ZN(n767) );
  NOR2_X1 U858 ( .A1(G1966), .A2(n806), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G2084), .A2(n755), .ZN(n775) );
  NOR2_X1 U860 ( .A1(n777), .A2(n775), .ZN(n756) );
  NAND2_X1 U861 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U862 ( .A(KEYINPUT30), .B(n757), .ZN(n758) );
  NOR2_X1 U863 ( .A1(G168), .A2(n758), .ZN(n761) );
  NOR2_X1 U864 ( .A1(G171), .A2(n759), .ZN(n760) );
  NOR2_X1 U865 ( .A1(n761), .A2(n760), .ZN(n764) );
  INV_X1 U866 ( .A(KEYINPUT31), .ZN(n762) );
  AND2_X1 U867 ( .A1(n773), .A2(n765), .ZN(n766) );
  OR2_X1 U868 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n779) );
  AND2_X1 U871 ( .A1(G8), .A2(n775), .ZN(n776) );
  NOR2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n798) );
  INV_X1 U874 ( .A(n806), .ZN(n780) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n946) );
  AND2_X1 U876 ( .A1(n780), .A2(n946), .ZN(n782) );
  AND2_X1 U877 ( .A1(n798), .A2(n782), .ZN(n781) );
  NAND2_X1 U878 ( .A1(n799), .A2(n781), .ZN(n788) );
  INV_X1 U879 ( .A(n782), .ZN(n786) );
  NOR2_X1 U880 ( .A1(G1976), .A2(G288), .ZN(n944) );
  NOR2_X1 U881 ( .A1(G1971), .A2(G303), .ZN(n783) );
  NOR2_X1 U882 ( .A1(n944), .A2(n783), .ZN(n784) );
  XNOR2_X1 U883 ( .A(n784), .B(KEYINPUT104), .ZN(n785) );
  OR2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n790) );
  XNOR2_X1 U886 ( .A(n790), .B(n789), .ZN(n792) );
  INV_X1 U887 ( .A(KEYINPUT33), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n944), .A2(KEYINPUT33), .ZN(n793) );
  NOR2_X1 U890 ( .A1(n793), .A2(n806), .ZN(n795) );
  XOR2_X1 U891 ( .A(G1981), .B(G305), .Z(n961) );
  NAND2_X1 U892 ( .A1(n796), .A2(n515), .ZN(n797) );
  XNOR2_X1 U893 ( .A(KEYINPUT105), .B(n797), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U896 ( .A1(G8), .A2(n800), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n806), .A2(n803), .ZN(n808) );
  NOR2_X1 U899 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XOR2_X1 U900 ( .A(n804), .B(KEYINPUT24), .Z(n805) );
  OR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n814) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n960) );
  NAND2_X1 U906 ( .A1(n960), .A2(n825), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n828) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n880), .ZN(n1006) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n852), .ZN(n1002) );
  NOR2_X1 U911 ( .A1(n815), .A2(n1002), .ZN(n818) );
  INV_X1 U912 ( .A(n816), .ZN(n817) );
  NOR2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n1006), .A2(n819), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n823), .A2(n883), .ZN(n1017) );
  NAND2_X1 U918 ( .A1(n824), .A2(n1017), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U924 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XNOR2_X1 U928 ( .A(G1348), .B(G2454), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n834), .B(G2430), .ZN(n835) );
  XNOR2_X1 U930 ( .A(n835), .B(G1341), .ZN(n841) );
  XOR2_X1 U931 ( .A(G2443), .B(G2427), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2438), .B(G2446), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n839) );
  XOR2_X1 U934 ( .A(G2451), .B(G2435), .Z(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n842), .A2(G14), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT106), .B(n843), .Z(G401) );
  INV_X1 U939 ( .A(n844), .ZN(G319) );
  NAND2_X1 U940 ( .A1(G124), .A2(n872), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U942 ( .A1(n870), .A2(G112), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G100), .A2(n614), .ZN(n849) );
  NAND2_X1 U945 ( .A1(G136), .A2(n867), .ZN(n848) );
  NAND2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U947 ( .A1(n851), .A2(n850), .ZN(G162) );
  XNOR2_X1 U948 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n852), .B(G162), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n864) );
  NAND2_X1 U951 ( .A1(G106), .A2(n614), .ZN(n856) );
  NAND2_X1 U952 ( .A1(G142), .A2(n867), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n857), .B(KEYINPUT45), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G130), .A2(n872), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U957 ( .A1(G118), .A2(n870), .ZN(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT111), .B(n860), .ZN(n861) );
  NOR2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U960 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U961 ( .A(G164), .B(n1001), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(n879) );
  NAND2_X1 U963 ( .A1(G103), .A2(n614), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G139), .A2(n867), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n878) );
  NAND2_X1 U966 ( .A1(n870), .A2(G115), .ZN(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT113), .B(n871), .ZN(n875) );
  NAND2_X1 U968 ( .A1(n872), .A2(G127), .ZN(n873) );
  XOR2_X1 U969 ( .A(KEYINPUT112), .B(n873), .Z(n874) );
  NOR2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U971 ( .A(n876), .B(KEYINPUT47), .ZN(n877) );
  NOR2_X1 U972 ( .A1(n878), .A2(n877), .ZN(n997) );
  XOR2_X1 U973 ( .A(n879), .B(n997), .Z(n882) );
  XOR2_X1 U974 ( .A(G160), .B(n880), .Z(n881) );
  XNOR2_X1 U975 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U976 ( .A(n884), .B(n883), .Z(n885) );
  NOR2_X1 U977 ( .A1(G37), .A2(n885), .ZN(G395) );
  XOR2_X1 U978 ( .A(n886), .B(G286), .Z(n888) );
  XNOR2_X1 U979 ( .A(n943), .B(n950), .ZN(n887) );
  XNOR2_X1 U980 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U981 ( .A(n889), .B(G171), .ZN(n890) );
  NOR2_X1 U982 ( .A1(G37), .A2(n890), .ZN(G397) );
  XOR2_X1 U983 ( .A(KEYINPUT108), .B(G2678), .Z(n892) );
  XNOR2_X1 U984 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n891) );
  XNOR2_X1 U985 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U986 ( .A(KEYINPUT42), .B(G2090), .Z(n894) );
  XNOR2_X1 U987 ( .A(G2067), .B(G2072), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U990 ( .A(G2096), .B(G2100), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U992 ( .A(G2084), .B(G2078), .Z(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(G227) );
  XNOR2_X1 U994 ( .A(G1981), .B(G2474), .ZN(n910) );
  XOR2_X1 U995 ( .A(G1976), .B(G1956), .Z(n902) );
  XNOR2_X1 U996 ( .A(G1966), .B(G1961), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U998 ( .A(G1971), .B(G1986), .Z(n904) );
  XNOR2_X1 U999 ( .A(G1996), .B(G1991), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1001 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1002 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(G229) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n911), .B(KEYINPUT114), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n913), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n914) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(G225) );
  XNOR2_X1 U1012 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(G325) );
  INV_X1 U1018 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1019 ( .A(G5), .B(n919), .ZN(n937) );
  XOR2_X1 U1020 ( .A(G1348), .B(KEYINPUT59), .Z(n920) );
  XNOR2_X1 U1021 ( .A(G4), .B(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G20), .B(G1956), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1341), .B(G19), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G1981), .B(G6), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT60), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(G1986), .B(G24), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G23), .B(G1976), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1032 ( .A(G1971), .B(KEYINPUT126), .Z(n930) );
  XNOR2_X1 U1033 ( .A(G22), .B(n930), .ZN(n931) );
  NAND2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(G21), .B(G1966), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1040 ( .A(KEYINPUT61), .B(n940), .Z(n941) );
  NOR2_X1 U1041 ( .A1(G16), .A2(n941), .ZN(n942) );
  XOR2_X1 U1042 ( .A(KEYINPUT127), .B(n942), .Z(n1026) );
  XOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .Z(n969) );
  XNOR2_X1 U1044 ( .A(G171), .B(G1961), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(n943), .B(G1348), .ZN(n949) );
  INV_X1 U1046 ( .A(n944), .ZN(n945) );
  NAND2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1048 ( .A(KEYINPUT124), .B(n947), .Z(n948) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n953) );
  XOR2_X1 U1050 ( .A(G1341), .B(n950), .Z(n951) );
  XNOR2_X1 U1051 ( .A(KEYINPUT125), .B(n951), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G166), .B(G1971), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(G1956), .B(KEYINPUT123), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(n956), .B(G299), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(n963), .B(KEYINPUT57), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n994) );
  XNOR2_X1 U1065 ( .A(G1991), .B(G25), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(G27), .B(n970), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G1996), .B(G32), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(G33), .B(G2072), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT120), .B(G2067), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(G26), .B(n975), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT121), .B(n978), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(G28), .A2(n981), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(n982), .B(KEYINPUT53), .ZN(n985) );
  XOR2_X1 U1078 ( .A(G2084), .B(G34), .Z(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT54), .B(n983), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G35), .B(G2090), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(KEYINPUT55), .B(n988), .ZN(n990) );
  INV_X1 U1084 ( .A(G29), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n991), .A2(G11), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT122), .B(n992), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n1024) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n995) );
  XNOR2_X1 U1090 ( .A(KEYINPUT118), .B(n995), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n997), .B(n996), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1000), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(G160), .B(G2084), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1007), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT119), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1019), .ZN(n1021) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(G29), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(n1027), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

