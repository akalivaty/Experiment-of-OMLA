//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(new_n191), .A3(G143), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n193), .B(G146), .C1(new_n189), .C2(KEYINPUT1), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n198), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n210), .B(KEYINPUT10), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT11), .B1(new_n212), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G134), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n213), .A2(new_n216), .B1(new_n212), .B2(G137), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(G101), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT78), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT78), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n219), .A2(new_n220), .A3(new_n223), .A4(G101), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT0), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n189), .A3(KEYINPUT64), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(KEYINPUT0), .B2(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n227), .B1(new_n233), .B2(new_n226), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n219), .A2(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n225), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n211), .A2(new_n218), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT76), .B(G140), .Z(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G227), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n240), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT75), .B(G110), .Z(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n206), .A2(new_n209), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n212), .A2(G137), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n214), .B1(G134), .B2(new_n215), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n212), .A2(KEYINPUT11), .A3(G137), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n257), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n251), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n251), .A2(KEYINPUT79), .A3(KEYINPUT12), .A4(new_n259), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n250), .A2(new_n266), .A3(new_n210), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n259), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n250), .B2(new_n210), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n247), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n218), .B1(new_n211), .B2(new_n238), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n246), .B1(new_n273), .B2(new_n239), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n187), .B(new_n188), .C1(new_n271), .C2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n187), .A2(new_n188), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n247), .A2(new_n272), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n262), .A3(new_n263), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n239), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT81), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n283), .A3(new_n239), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n279), .B1(new_n285), .B2(new_n245), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n278), .B1(new_n286), .B2(G469), .ZN(new_n287));
  INV_X1    g101(.A(G221), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT9), .B(G234), .Z(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n188), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT82), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n280), .A2(new_n283), .A3(new_n239), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n283), .B1(new_n280), .B2(new_n239), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n245), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n279), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(G469), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n280), .A2(new_n246), .A3(new_n239), .ZN(new_n297));
  INV_X1    g111(.A(new_n239), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n245), .B1(new_n298), .B2(new_n272), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n276), .B1(new_n300), .B2(new_n187), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n303));
  INV_X1    g117(.A(new_n290), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n307), .A2(KEYINPUT16), .A3(G140), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT16), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n191), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n309), .B(G146), .C1(new_n313), .C2(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n308), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n321), .A2(new_n317), .A3(G146), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT24), .B(G110), .Z(new_n324));
  XNOR2_X1  g138(.A(G119), .B(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT23), .B1(new_n189), .B2(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n189), .A2(G119), .ZN(new_n328));
  MUX2_X1   g142(.A(KEYINPUT23), .B(new_n327), .S(new_n328), .Z(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G110), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n319), .A2(new_n323), .A3(new_n326), .A4(new_n330), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n329), .A2(G110), .B1(new_n325), .B2(new_n324), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n318), .C1(G146), .C2(new_n313), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G137), .ZN(new_n335));
  INV_X1    g149(.A(G234), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n288), .A2(new_n336), .A3(G953), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n335), .B(new_n337), .Z(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n333), .A3(new_n338), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n188), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT25), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT72), .B(G217), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(G234), .B2(new_n188), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(KEYINPUT25), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n344), .A2(KEYINPUT25), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n342), .A2(new_n188), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n348), .A2(G902), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n215), .B2(G134), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n215), .A2(G134), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n212), .A2(KEYINPUT65), .A3(G137), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G131), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n198), .A3(new_n258), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n198), .A2(new_n361), .A3(new_n258), .A4(KEYINPUT66), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n364), .B(new_n365), .C1(new_n218), .C2(new_n234), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT30), .B(new_n362), .C1(new_n218), .C2(new_n234), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n370));
  INV_X1    g184(.A(G113), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT67), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT67), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(KEYINPUT2), .B2(G113), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n372), .A2(new_n374), .B1(KEYINPUT2), .B2(G113), .ZN(new_n375));
  XNOR2_X1  g189(.A(G116), .B(G119), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n369), .A3(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n375), .A2(new_n376), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n362), .C1(new_n218), .C2(new_n234), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT26), .B(G101), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n241), .A3(G210), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n383), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n378), .A2(new_n382), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT31), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n378), .A2(KEYINPUT31), .A3(new_n382), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n234), .B1(new_n256), .B2(new_n258), .ZN(new_n397));
  INV_X1    g211(.A(new_n362), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n397), .A2(new_n398), .A3(new_n377), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT28), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n377), .B2(new_n366), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT69), .ZN(new_n404));
  INV_X1    g218(.A(new_n390), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n388), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n389), .A2(KEYINPUT69), .A3(new_n390), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(G472), .A2(G902), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT32), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n394), .A2(new_n395), .B1(new_n403), .B2(new_n408), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT32), .ZN(new_n414));
  INV_X1    g228(.A(new_n411), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n377), .B1(new_n397), .B2(new_n398), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT71), .A3(new_n382), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT71), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n377), .C1(new_n397), .C2(new_n398), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(KEYINPUT28), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n400), .A3(new_n391), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n423), .A2(KEYINPUT29), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n406), .A2(new_n407), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n400), .B(new_n426), .C1(new_n401), .C2(new_n402), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n397), .A2(new_n398), .A3(new_n367), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n367), .B2(new_n366), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n399), .B1(new_n429), .B2(new_n377), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n427), .B1(new_n430), .B2(new_n391), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n188), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G472), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n355), .B1(new_n417), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n225), .A2(new_n377), .A3(new_n237), .ZN(new_n439));
  INV_X1    g253(.A(new_n249), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n375), .A2(new_n376), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n442));
  INV_X1    g256(.A(G116), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G119), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT5), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n371), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n440), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n438), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n450), .B(new_n437), .C1(new_n439), .C2(new_n448), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n439), .A2(new_n450), .A3(new_n448), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n235), .A2(G125), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n198), .A2(new_n307), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G224), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n456), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n457), .B2(new_n458), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n450), .B(KEYINPUT8), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n446), .A2(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n442), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n446), .A2(KEYINPUT85), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n441), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n469), .B2(new_n440), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n441), .A2(new_n249), .A3(new_n447), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n464), .A2(KEYINPUT7), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT86), .B(KEYINPUT7), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(new_n461), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(new_n454), .C1(new_n459), .C2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n475), .A2(new_n188), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n449), .A2(new_n451), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n437), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n449), .A2(new_n451), .A3(new_n438), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n454), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n481));
  INV_X1    g295(.A(new_n462), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n463), .A2(new_n476), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n463), .A2(new_n476), .A3(new_n485), .A4(new_n483), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n436), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n384), .A2(new_n241), .A3(G214), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n193), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G131), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n490), .B(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n257), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n493), .A2(new_n257), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT17), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n318), .A2(new_n317), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n321), .A2(G146), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n496), .B(new_n498), .C1(new_n501), .C2(new_n322), .ZN(new_n502));
  XNOR2_X1  g316(.A(G113), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n199), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT18), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n493), .B1(new_n505), .B2(new_n257), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n320), .B(new_n191), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n507), .C1(new_n505), .C2(new_n492), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n502), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n320), .B(KEYINPUT19), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n191), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n491), .A2(G131), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n318), .C1(new_n497), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n508), .ZN(new_n514));
  INV_X1    g328(.A(new_n504), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT20), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT88), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n517), .A2(new_n522), .A3(new_n518), .A4(new_n519), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n519), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n509), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n504), .B1(new_n502), .B2(new_n508), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n188), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G475), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n346), .A2(new_n289), .A3(new_n241), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n443), .A2(G122), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n536));
  INV_X1    g350(.A(G122), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(G116), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n443), .A2(KEYINPUT89), .A3(G122), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT90), .B(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n543), .B1(new_n544), .B2(new_n534), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n538), .A2(new_n539), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n542), .B(new_n545), .C1(KEYINPUT14), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G107), .ZN(new_n548));
  XNOR2_X1  g362(.A(G128), .B(G143), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(new_n212), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n202), .A3(new_n535), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(KEYINPUT13), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n193), .A2(G128), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n555), .B(G134), .C1(KEYINPUT13), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n212), .ZN(new_n558));
  INV_X1    g372(.A(new_n551), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n202), .B1(new_n546), .B2(new_n535), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(KEYINPUT91), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n552), .B1(new_n547), .B2(G107), .ZN(new_n564));
  INV_X1    g378(.A(new_n561), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n533), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n533), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(KEYINPUT91), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n188), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n188), .B(new_n579), .C1(new_n567), .C2(new_n570), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n241), .A2(G952), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n336), .B2(new_n384), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT21), .B(G898), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT93), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n188), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n532), .A2(new_n581), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n489), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n306), .A2(new_n434), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT94), .B(G101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G3));
  INV_X1    g408(.A(new_n355), .ZN(new_n595));
  OAI21_X1  g409(.A(G472), .B1(new_n413), .B2(G902), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n410), .A2(new_n411), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n306), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n291), .B2(new_n305), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT95), .A3(new_n595), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n589), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n567), .B2(new_n570), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n572), .A2(G902), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n568), .A2(KEYINPUT96), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n569), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n569), .A2(new_n610), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n571), .A2(new_n572), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n616), .A2(new_n532), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n489), .A2(new_n606), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n489), .A2(KEYINPUT97), .A3(new_n606), .A4(new_n617), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n605), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n525), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n517), .A2(new_n519), .A3(new_n625), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n526), .A2(new_n626), .B1(new_n530), .B2(G475), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n581), .A2(new_n606), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n581), .A2(KEYINPUT98), .A3(new_n606), .A4(new_n627), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n630), .A2(new_n489), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n605), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n334), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n353), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n352), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n603), .A2(new_n591), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(new_n489), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n584), .B1(new_n588), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n581), .A2(new_n627), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n639), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n417), .B2(new_n433), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n306), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  NAND2_X1  g466(.A1(new_n487), .A2(new_n488), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n419), .A2(new_n421), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n430), .A2(new_n391), .B1(new_n657), .B2(new_n408), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n658), .B2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n417), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n532), .A2(new_n581), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n649), .A2(new_n662), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n655), .A2(new_n661), .A3(new_n436), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n645), .B(KEYINPUT39), .Z(new_n665));
  AOI21_X1  g479(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n666));
  AOI211_X1 g480(.A(KEYINPUT82), .B(new_n290), .C1(new_n296), .C2(new_n301), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT100), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n665), .C1(new_n666), .C2(new_n667), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n669), .A2(KEYINPUT40), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT40), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n664), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  AND3_X1   g489(.A1(new_n616), .A2(new_n532), .A3(new_n646), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n489), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n489), .A2(new_n676), .A3(KEYINPUT101), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n306), .A3(new_n650), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NAND3_X1  g496(.A1(new_n410), .A2(KEYINPUT32), .A3(new_n411), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n433), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n300), .A2(new_n187), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n686), .A2(new_n304), .A3(new_n275), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n685), .A2(new_n595), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n620), .A2(new_n621), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND2_X1  g505(.A1(new_n632), .A2(new_n688), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  AND3_X1   g507(.A1(new_n685), .A2(new_n639), .A3(new_n687), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(KEYINPUT102), .A3(new_n591), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n685), .A2(new_n639), .A3(new_n687), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n489), .A2(new_n590), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  NAND2_X1  g515(.A1(new_n422), .A2(new_n400), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n408), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n415), .B1(new_n396), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n596), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(KEYINPUT103), .B(G472), .C1(new_n413), .C2(G902), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n704), .B(new_n355), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n489), .A2(new_n662), .A3(new_n687), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n606), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  AOI211_X1 g525(.A(new_n704), .B(new_n649), .C1(new_n706), .C2(new_n707), .ZN(new_n712));
  INV_X1    g526(.A(new_n687), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n677), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n412), .B2(new_n416), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT104), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n433), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n595), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n487), .A2(new_n435), .A3(new_n488), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n287), .A3(new_n290), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n676), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT42), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n434), .A2(new_n723), .A3(new_n726), .A4(new_n676), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n257), .ZN(G33));
  OR2_X1    g543(.A1(new_n647), .A2(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n647), .A2(KEYINPUT105), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n434), .A2(new_n723), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  NAND3_X1  g547(.A1(new_n294), .A2(KEYINPUT45), .A3(new_n295), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n246), .B1(new_n282), .B2(new_n284), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n279), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n294), .A2(KEYINPUT106), .A3(KEYINPUT45), .A4(new_n295), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(G469), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n277), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n277), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n275), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n304), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n532), .A2(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n532), .A2(KEYINPUT107), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n616), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT43), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n532), .A2(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n616), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n598), .A3(new_n639), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n722), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n747), .A2(new_n756), .A3(new_n665), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  NOR3_X1   g573(.A1(new_n685), .A2(new_n722), .A3(new_n595), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n745), .A2(new_n275), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT46), .B1(new_n741), .B2(new_n277), .ZN(new_n762));
  OAI211_X1 g576(.A(KEYINPUT47), .B(new_n304), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT47), .B1(new_n746), .B2(new_n304), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n676), .B(new_n760), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  AND4_X1   g581(.A1(new_n584), .A2(new_n751), .A3(new_n708), .A4(new_n753), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n687), .ZN(new_n769));
  INV_X1    g583(.A(new_n655), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n769), .A2(new_n435), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT50), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n764), .A2(new_n765), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n686), .A2(new_n275), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n304), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n722), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n768), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n713), .A2(new_n722), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n584), .A2(new_n751), .A3(new_n753), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n712), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n661), .A2(new_n780), .A3(new_n595), .A4(new_n584), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n783), .A2(new_n532), .A3(new_n616), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n779), .A2(KEYINPUT109), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n782), .A2(new_n786), .A3(KEYINPUT51), .A4(new_n784), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n689), .A2(new_n710), .A3(new_n692), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT102), .B1(new_n694), .B2(new_n591), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n697), .A2(new_n698), .A3(new_n696), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n489), .A2(new_n662), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n589), .A3(new_n713), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n799), .A2(new_n708), .B1(new_n632), .B2(new_n688), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n700), .A3(KEYINPUT108), .A4(new_n689), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n643), .A2(new_n589), .ZN(new_n803));
  INV_X1    g617(.A(new_n617), .ZN(new_n804));
  INV_X1    g618(.A(new_n581), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n805), .B2(new_n532), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n602), .A2(new_n604), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n640), .A2(new_n592), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n725), .A2(new_n727), .A3(new_n732), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n712), .A2(new_n676), .A3(new_n723), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n627), .A2(new_n646), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n306), .A2(new_n650), .A3(new_n805), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n814), .B2(new_n722), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n681), .A2(new_n715), .A3(new_n651), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n643), .A2(new_n663), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n287), .A2(new_n290), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n646), .A4(new_n660), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n681), .A3(new_n715), .A4(new_n651), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n791), .B1(new_n810), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n793), .A2(new_n796), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n808), .A4(new_n807), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n823), .B(new_n818), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n816), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n807), .A2(new_n808), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n797), .B2(new_n801), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n816), .A3(new_n830), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n791), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n833), .B1(new_n837), .B2(KEYINPUT54), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n781), .A2(new_n595), .A3(new_n720), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT48), .Z(new_n840));
  OAI221_X1 g654(.A(new_n582), .B1(new_n804), .B2(new_n783), .C1(new_n769), .C2(new_n643), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT110), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n790), .A2(new_n844), .B1(G952), .B2(G953), .ZN(new_n845));
  INV_X1    g659(.A(new_n750), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n595), .C1(KEYINPUT49), .C2(new_n775), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n770), .B(new_n847), .C1(KEYINPUT49), .C2(new_n775), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n304), .A3(new_n435), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n845), .B1(new_n660), .B2(new_n849), .ZN(G75));
  NOR2_X1   g664(.A1(new_n241), .A2(G952), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT114), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n825), .A2(new_n828), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n836), .B2(new_n791), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n188), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT56), .B1(new_n856), .B2(G210), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n480), .B(KEYINPUT111), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT55), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n462), .B(KEYINPUT112), .Z(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(KEYINPUT113), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n853), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n857), .B2(new_n863), .ZN(G51));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n855), .A2(new_n188), .A3(new_n741), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n855), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n277), .A2(KEYINPUT57), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n276), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n297), .A2(new_n299), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n866), .B1(new_n877), .B2(new_n851), .ZN(new_n878));
  INV_X1    g692(.A(new_n851), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n276), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n880), .A2(new_n872), .B1(new_n299), .B2(new_n297), .ZN(new_n881));
  OAI211_X1 g695(.A(KEYINPUT115), .B(new_n879), .C1(new_n881), .C2(new_n867), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(G54));
  NAND3_X1  g697(.A1(new_n856), .A2(KEYINPUT58), .A3(G475), .ZN(new_n884));
  INV_X1    g698(.A(new_n517), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n884), .A2(KEYINPUT116), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n851), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT116), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G60));
  AND2_X1   g703(.A1(new_n608), .A2(new_n613), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n572), .A2(new_n188), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n891), .B(new_n892), .Z(new_n893));
  NAND3_X1  g707(.A1(new_n871), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n893), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n838), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n853), .B(new_n894), .C1(new_n896), .C2(new_n890), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(G63));
  INV_X1    g712(.A(new_n342), .ZN(new_n899));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT60), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n855), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n826), .B2(new_n831), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n637), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n902), .A2(new_n904), .A3(KEYINPUT61), .A4(new_n853), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n902), .B2(new_n853), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n908), .B(new_n853), .C1(new_n903), .C2(new_n342), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n906), .B(new_n907), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n853), .B1(new_n903), .B2(new_n342), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT118), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n910), .A3(new_n904), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n906), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n905), .B1(new_n913), .B2(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n587), .B2(new_n460), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n835), .A2(G953), .B1(KEYINPUT120), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(KEYINPUT120), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n858), .B1(G898), .B2(new_n241), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n921), .B(new_n922), .Z(G69));
  AOI21_X1  g737(.A(new_n241), .B1(G227), .B2(G900), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT124), .Z(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n655), .A2(new_n663), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n435), .A3(new_n660), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT40), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n670), .B1(new_n306), .B2(new_n665), .ZN(new_n932));
  INV_X1    g746(.A(new_n671), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n669), .A2(KEYINPUT40), .A3(new_n671), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n930), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n681), .A2(new_n715), .A3(new_n651), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT62), .B1(new_n674), .B2(new_n817), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n932), .A2(new_n933), .A3(new_n722), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n434), .A3(new_n806), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n766), .A2(new_n758), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n928), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n766), .A2(new_n758), .A3(new_n943), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n937), .B1(new_n936), .B2(new_n938), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n674), .A2(KEYINPUT62), .A3(new_n817), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT122), .ZN(new_n950));
  AOI21_X1  g764(.A(G953), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n510), .B(KEYINPUT121), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n429), .B(new_n952), .Z(new_n953));
  OAI21_X1  g767(.A(new_n927), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT122), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT122), .B1(new_n946), .B2(new_n949), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n241), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n953), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(KEYINPUT123), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n961));
  INV_X1    g775(.A(new_n811), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n758), .A2(new_n766), .A3(new_n962), .A4(new_n817), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n747), .A2(new_n665), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n964), .A2(new_n798), .A3(new_n721), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT125), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n766), .A2(new_n758), .A3(new_n962), .A4(new_n817), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n965), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n241), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n241), .A2(G900), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n953), .ZN(new_n975));
  AND4_X1   g789(.A1(new_n926), .A2(new_n960), .A3(new_n961), .A4(new_n975), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n954), .A2(new_n959), .B1(new_n974), .B2(new_n953), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n926), .B1(new_n977), .B2(new_n961), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n976), .A2(new_n978), .ZN(G72));
  INV_X1    g793(.A(new_n430), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n391), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n391), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n837), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT127), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n955), .A2(new_n956), .A3(new_n810), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n391), .B(new_n980), .C1(new_n989), .C2(new_n984), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n967), .A2(new_n970), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n983), .B1(new_n991), .B2(new_n810), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n851), .B1(new_n992), .B2(new_n981), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n988), .A2(new_n990), .A3(new_n993), .ZN(G57));
endmodule


