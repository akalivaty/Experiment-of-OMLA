//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(new_n459), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n472), .B(new_n460), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(new_n467), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT68), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n475), .A2(KEYINPUT68), .A3(new_n476), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  NAND4_X1  g057(.A1(new_n464), .A2(G2105), .A3(new_n465), .A4(new_n467), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT71), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n468), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G136), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n465), .A3(new_n467), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n475), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n459), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n483), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n500), .A2(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n506), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT74), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(new_n519), .A3(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n509), .A2(new_n511), .B1(new_n508), .B2(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n510), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n524), .A2(G88), .B1(G50), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n520), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND2_X1   g105(.A1(new_n524), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n527), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n527), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n523), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(G64), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR3_X1    g119(.A1(new_n540), .A2(new_n544), .A3(KEYINPUT75), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT75), .B1(new_n540), .B2(new_n544), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n527), .A2(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n523), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n541), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n514), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n557), .A2(KEYINPUT76), .A3(G651), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n551), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n521), .A2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n521), .A2(G91), .A3(new_n522), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n522), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n527), .A2(new_n574), .A3(G53), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n569), .A2(new_n570), .A3(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  OAI21_X1  g154(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI221_X1 g157(.A(new_n580), .B1(new_n581), .B2(new_n571), .C1(new_n582), .C2(new_n523), .ZN(G288));
  NAND2_X1  g158(.A1(new_n527), .A2(G48), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n541), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n521), .A2(G86), .A3(new_n522), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n514), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(KEYINPUT78), .A3(G651), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n527), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n523), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n521), .A2(G92), .A3(new_n522), .A4(new_n604), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n607), .A2(new_n608), .B1(G54), .B2(new_n527), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n514), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g189(.A(KEYINPUT80), .B(new_n610), .C1(new_n514), .C2(new_n611), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n614), .A2(G651), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n603), .B1(new_n619), .B2(new_n602), .ZN(G284));
  AOI21_X1  g195(.A(new_n603), .B1(new_n619), .B2(new_n602), .ZN(G321));
  NOR2_X1   g196(.A1(G286), .A2(new_n602), .ZN(new_n622));
  XNOR2_X1  g197(.A(G299), .B(KEYINPUT82), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n602), .ZN(G297));
  AOI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n602), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NOR2_X1   g202(.A1(new_n560), .A2(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n619), .A2(new_n626), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n459), .A2(G2104), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n475), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n634), .B(new_n635), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2100), .Z(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n483), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G135), .B2(new_n490), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n638), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n650), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n664), .A2(new_n649), .A3(new_n660), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  OAI21_X1  g242(.A(KEYINPUT86), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(new_n667), .ZN(new_n670));
  NAND4_X1  g245(.A1(new_n663), .A2(new_n665), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G14), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n667), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(G401));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  OR3_X1    g254(.A1(new_n678), .A2(KEYINPUT87), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT87), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(new_n676), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n677), .B(KEYINPUT17), .Z(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n676), .A3(new_n677), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT18), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n679), .A3(new_n682), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n694), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n694), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR3_X1    g279(.A1(new_n700), .A2(new_n704), .A3(KEYINPUT88), .ZN(new_n705));
  OAI21_X1  g280(.A(KEYINPUT88), .B1(new_n700), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n705), .B2(new_n706), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n691), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(new_n691), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n713), .A3(new_n708), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n711), .B2(new_n714), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(G229));
  NOR2_X1   g293(.A1(G29), .A2(G35), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G162), .B2(G29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2090), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT100), .Z(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G33), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT95), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT25), .ZN(new_n729));
  NAND2_X1  g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  INV_X1    g305(.A(G127), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n475), .B2(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n728), .A2(new_n729), .B1(G2105), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n490), .A2(G139), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n725), .B1(new_n736), .B2(new_n724), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2072), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G164), .A2(new_n724), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G27), .B2(new_n724), .ZN(new_n745));
  INV_X1    g320(.A(G2078), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n743), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n644), .B2(new_n724), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n643), .A2(KEYINPUT98), .A3(G29), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  OR3_X1    g328(.A1(new_n753), .A2(KEYINPUT99), .A3(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT99), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n751), .A2(new_n752), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n738), .A2(new_n749), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n739), .A2(G4), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n619), .B2(new_n739), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(G1348), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G160), .A2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G34), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(new_n724), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT96), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2084), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n760), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n764), .B2(new_n762), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n721), .A2(G2090), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT89), .B(G16), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G19), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n560), .B2(new_n776), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT94), .B(G1341), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G5), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G171), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G129), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n483), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT26), .Z(new_n789));
  INV_X1    g364(.A(G105), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n633), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n490), .B2(G141), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n724), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n724), .B2(G32), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n775), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n570), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n541), .B1(new_n566), .B2(new_n567), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n804), .B2(new_n739), .ZN(new_n805));
  INV_X1    g380(.A(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n724), .A2(G26), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT28), .ZN(new_n809));
  INV_X1    g384(.A(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n459), .A2(G116), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n483), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G140), .B2(new_n490), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(new_n724), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n796), .B2(new_n797), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n784), .A2(new_n798), .A3(new_n807), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n774), .A2(new_n780), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n723), .A2(new_n773), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(KEYINPUT92), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n776), .A2(G24), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G290), .B2(new_n775), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT90), .B(G1986), .Z(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n724), .A2(G25), .ZN(new_n828));
  OR2_X1    g403(.A1(G95), .A2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n830));
  INV_X1    g405(.A(G119), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n483), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G131), .B2(new_n490), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n828), .B1(new_n833), .B2(new_n724), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G1991), .Z(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n825), .B2(new_n826), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n776), .A2(G22), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n776), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G1971), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n739), .A2(G23), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n523), .A2(new_n582), .B1(new_n581), .B2(new_n571), .ZN(new_n845));
  INV_X1    g420(.A(new_n580), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n844), .B1(new_n847), .B2(new_n739), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT33), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1976), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n739), .A2(G6), .ZN(new_n851));
  INV_X1    g426(.A(G305), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n739), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT32), .B(G1981), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n843), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT91), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT34), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n840), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(KEYINPUT34), .A3(new_n859), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n823), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n823), .A3(new_n863), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n820), .B1(new_n865), .B2(new_n866), .ZN(G311));
  INV_X1    g442(.A(new_n820), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n864), .ZN(G150));
  NAND3_X1  g445(.A1(new_n512), .A2(G67), .A3(new_n513), .ZN(new_n871));
  NAND2_X1  g446(.A1(G80), .A2(G543), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G651), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n512), .A2(G93), .A3(new_n513), .A4(new_n522), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(G55), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n527), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n876), .B1(new_n875), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G860), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n619), .A2(G559), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n884), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(KEYINPUT105), .B(new_n874), .C1(new_n879), .C2(new_n880), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n559), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n880), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n892), .A2(new_n893), .B1(G651), .B2(new_n873), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n557), .A2(G651), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n550), .B1(new_n895), .B2(new_n552), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n894), .A2(new_n896), .A3(KEYINPUT105), .A4(new_n558), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n887), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n900));
  AOI21_X1  g475(.A(G860), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n900), .B2(new_n899), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n883), .B1(new_n903), .B2(new_n904), .ZN(G145));
  OR2_X1    g480(.A1(G162), .A2(G160), .ZN(new_n906));
  NAND2_X1  g481(.A1(G162), .A2(G160), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n643), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n643), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n636), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n833), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n490), .A2(G142), .ZN(new_n915));
  INV_X1    g490(.A(G130), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n459), .A2(G118), .ZN(new_n917));
  OAI21_X1  g492(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n918));
  OAI221_X1 g493(.A(new_n915), .B1(new_n916), .B2(new_n483), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n914), .A2(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n912), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n914), .A2(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n636), .A3(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n814), .B(G164), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n736), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n736), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n794), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n793), .B1(new_n934), .B2(new_n930), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n927), .A2(new_n928), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n933), .A3(new_n923), .A4(new_n925), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n926), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n911), .A2(new_n936), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n910), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n908), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n937), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g522(.A(new_n629), .B(new_n898), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n617), .A2(KEYINPUT109), .A3(G299), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT109), .B1(new_n802), .B2(new_n803), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n569), .A2(new_n951), .A3(new_n570), .A4(new_n576), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n950), .A2(new_n616), .A3(new_n609), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n949), .B2(new_n953), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n948), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n949), .A2(new_n953), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT110), .Z(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n948), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n852), .A2(G303), .ZN(new_n965));
  NOR2_X1   g540(.A1(G166), .A2(G305), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(G288), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G290), .B(new_n847), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n970), .A2(new_n965), .A3(new_n966), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n964), .A2(KEYINPUT112), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n959), .A2(new_n975), .A3(new_n963), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n959), .B2(new_n963), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n973), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G868), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G868), .B2(new_n894), .ZN(G295));
  OAI21_X1  g556(.A(new_n980), .B1(G868), .B2(new_n894), .ZN(G331));
  AND3_X1   g557(.A1(new_n891), .A2(G171), .A3(new_n897), .ZN(new_n983));
  AOI21_X1  g558(.A(G171), .B1(new_n891), .B2(new_n897), .ZN(new_n984));
  OAI21_X1  g559(.A(G286), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n898), .A2(G301), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n891), .A2(new_n897), .A3(G171), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(G168), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n960), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n958), .B1(new_n985), .B2(new_n988), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n969), .A2(new_n971), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n961), .A2(new_n988), .A3(new_n985), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n960), .A2(KEYINPUT41), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n956), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n983), .A2(new_n984), .A3(G286), .ZN(new_n999));
  AOI21_X1  g574(.A(G168), .B1(new_n986), .B2(new_n987), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n997), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n1001), .A3(new_n972), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n994), .A2(new_n995), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n958), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n999), .B2(new_n1000), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n993), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G37), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n993), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(KEYINPUT114), .A3(new_n1006), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1003), .B1(new_n1014), .B2(new_n995), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT44), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n995), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n994), .A2(new_n1002), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1016), .A2(new_n1021), .ZN(G397));
  INV_X1    g597(.A(new_n473), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n465), .A2(new_n467), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(G137), .A3(new_n459), .A4(new_n464), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n472), .B1(new_n1025), .B2(new_n460), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n481), .B(G40), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n500), .B2(new_n504), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT115), .B(KEYINPUT45), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1996), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n793), .B(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n814), .B(G2067), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n833), .A2(new_n835), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n833), .A2(new_n835), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(G290), .B(G1986), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n587), .A2(new_n590), .A3(new_n1042), .A4(new_n591), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n586), .B2(new_n588), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(KEYINPUT120), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(KEYINPUT120), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1044), .A2(KEYINPUT120), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(KEYINPUT49), .A3(new_n1046), .A4(new_n1043), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  OAI221_X1 g630(.A(G8), .B1(new_n1055), .B2(G288), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G288), .A2(new_n1055), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g636(.A(KEYINPUT118), .B(KEYINPUT52), .C1(G288), .C2(new_n1055), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1056), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT119), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1066), .A2(new_n1056), .A3(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1054), .B(new_n1057), .C1(new_n1065), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT45), .B(new_n1028), .C1(new_n500), .C2(new_n504), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(new_n474), .A3(G40), .A4(new_n481), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1029), .A2(new_n1075), .A3(new_n1030), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1027), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n1028), .C1(new_n500), .C2(new_n504), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1078), .A2(G1971), .B1(new_n1083), .B2(G2090), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1072), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1069), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(G8), .A3(new_n1072), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1084), .A2(new_n1072), .A3(new_n1089), .A4(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1086), .A2(new_n1091), .A3(KEYINPUT125), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT125), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1073), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1027), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1077), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1029), .A2(new_n1075), .A3(new_n1030), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n804), .B(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n806), .B1(new_n1103), .B2(new_n1027), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1095), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OR3_X1    g684(.A1(new_n1105), .A2(new_n1106), .A3(new_n1095), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT123), .B(new_n1095), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1111));
  NAND2_X1  g686(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1049), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1078), .B2(new_n1033), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1113), .B1(new_n1116), .B2(new_n559), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G1996), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n560), .B(new_n1112), .C1(new_n1119), .C2(new_n1115), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n619), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n1103), .B2(new_n1027), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1079), .A2(new_n1125), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1126), .A3(new_n763), .ZN(new_n1127));
  INV_X1    g702(.A(G2067), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1049), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1127), .A2(KEYINPUT60), .A3(new_n619), .A4(new_n1129), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1106), .B1(new_n1130), .B2(new_n619), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1122), .A2(new_n1135), .B1(new_n1136), .B2(new_n1105), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1118), .B2(G2078), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1124), .A2(new_n1126), .A3(new_n783), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1097), .A2(KEYINPUT53), .A3(new_n746), .A4(new_n1031), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(G171), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT45), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1029), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1027), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(KEYINPUT53), .A3(new_n746), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1139), .A2(G301), .A3(new_n1140), .A4(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1143), .A2(KEYINPUT54), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n742), .B1(new_n1146), .B2(new_n1027), .ZN(new_n1152));
  INV_X1    g727(.A(G2084), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1079), .A2(new_n1153), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1151), .B(G8), .C1(new_n1155), .C2(G286), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G168), .A2(new_n1050), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1158), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT124), .B(new_n1160), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1156), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1151), .B(new_n1158), .C1(new_n1155), .C2(G8), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1139), .A2(new_n1148), .A3(new_n1140), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(G171), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1139), .A2(G301), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT54), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1150), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1137), .A2(new_n1169), .ZN(new_n1170));
  OR3_X1    g745(.A1(new_n1162), .A2(KEYINPUT62), .A3(new_n1163), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT62), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(G171), .A3(new_n1165), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1094), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1091), .A2(new_n1069), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1054), .A2(new_n1055), .A3(new_n847), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1043), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1175), .B1(new_n1051), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1050), .B(G286), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1086), .A2(new_n1091), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1178), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1040), .B1(new_n1174), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1035), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1032), .B1(new_n1186), .B2(new_n793), .ZN(new_n1187));
  NOR4_X1   g762(.A1(new_n1027), .A2(new_n1031), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT46), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1189), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1187), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT47), .ZN(new_n1192));
  NOR2_X1   g767(.A1(G290), .A2(G1986), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1032), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1038), .A2(new_n1032), .B1(KEYINPUT48), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(KEYINPUT48), .B2(new_n1195), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n814), .A2(new_n1128), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1036), .B(KEYINPUT126), .Z(new_n1200));
  OAI21_X1  g775(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1032), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1192), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1185), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(G319), .ZN(new_n1206));
  OR2_X1    g780(.A1(G227), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n672), .B2(new_n674), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1208), .B1(new_n716), .B2(new_n717), .ZN(new_n1209));
  AOI21_X1  g783(.A(new_n1209), .B1(new_n941), .B2(new_n945), .ZN(new_n1210));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n1015), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1011), .B1(new_n990), .B2(new_n991), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1212), .A2(new_n1013), .A3(new_n972), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n995), .B1(new_n1213), .B2(new_n994), .ZN(new_n1214));
  AND4_X1   g788(.A1(new_n1008), .A2(new_n1002), .A3(new_n995), .A4(new_n1007), .ZN(new_n1215));
  OAI211_X1 g789(.A(KEYINPUT127), .B(new_n1210), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  INV_X1    g790(.A(new_n1216), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1211), .A2(new_n1217), .ZN(G308));
  NAND2_X1  g792(.A1(new_n1015), .A2(new_n1210), .ZN(G225));
endmodule


