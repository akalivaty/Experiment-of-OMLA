//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n203), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n213), .B1(KEYINPUT1), .B2(new_n222), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n222), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n227), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT70), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(new_n226), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT64), .B(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(KEYINPUT70), .A3(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G77), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n262), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n255), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT79), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G68), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT12), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n267), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n253), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n207), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G68), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(KEYINPUT11), .B2(new_n264), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n265), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n265), .A2(new_n276), .A3(KEYINPUT80), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n236), .A2(G1698), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n282), .B1(G226), .B2(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT76), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n228), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT76), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(new_n292), .A3(new_n286), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n227), .B1(new_n298), .B2(new_n289), .ZN(new_n299));
  NAND3_X1  g0099(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G238), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n289), .A2(new_n298), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(new_n228), .A3(new_n300), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G274), .A3(new_n297), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n308));
  NAND3_X1  g0108(.A1(new_n294), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT78), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n294), .A2(new_n307), .ZN(new_n312));
  INV_X1    g0112(.A(new_n308), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n294), .A2(new_n307), .A3(KEYINPUT78), .A4(new_n308), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n293), .A2(new_n291), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n306), .B1(new_n319), .B2(new_n288), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT13), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n309), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n281), .A2(new_n317), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n316), .A2(new_n330), .A3(G169), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n281), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G222), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(G1698), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT68), .B(G223), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n339), .B1(new_n340), .B2(new_n337), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n291), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n301), .A2(G226), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(new_n305), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n323), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n344), .B2(new_n346), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n201), .B1(new_n207), .B2(G20), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n255), .A2(new_n267), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n271), .A2(new_n201), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n258), .A2(new_n260), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT71), .ZN(new_n359));
  NOR3_X1   g0159(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(new_n208), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n204), .A2(KEYINPUT71), .A3(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n262), .A2(G150), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n255), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n355), .B1(KEYINPUT72), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n358), .A2(new_n364), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n252), .A2(new_n227), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n254), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n366), .A2(new_n367), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n367), .B1(new_n366), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n351), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n379));
  OR2_X1    g0179(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n366), .A2(new_n375), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT9), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n366), .A2(new_n367), .A3(new_n375), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n385), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n351), .ZN(new_n386));
  INV_X1    g0186(.A(new_n382), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n347), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(G179), .B2(new_n347), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n381), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n372), .A2(new_n271), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n356), .B1(new_n207), .B2(G20), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(new_n271), .B2(new_n356), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n335), .A2(new_n223), .A3(new_n225), .A4(new_n336), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n283), .A2(new_n284), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n208), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(G68), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT81), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G58), .A3(G68), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n406), .A3(new_n230), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(G20), .B1(G159), .B2(new_n262), .ZN(new_n408));
  AOI211_X1 g0208(.A(KEYINPUT82), .B(KEYINPUT16), .C1(new_n402), .C2(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n283), .A2(new_n284), .A3(G20), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n410), .B2(new_n400), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n408), .B(KEYINPUT16), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n253), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(new_n408), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT82), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n396), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(G223), .B(new_n338), .C1(new_n283), .C2(new_n284), .ZN(new_n421));
  OAI211_X1 g0221(.A(G226), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n424), .A2(new_n291), .ZN(new_n425));
  INV_X1    g0225(.A(new_n297), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n304), .A2(new_n426), .A3(G232), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n305), .A2(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n425), .A2(new_n328), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n305), .A2(new_n427), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n424), .A2(new_n291), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n388), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n420), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT82), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n400), .B1(new_n399), .B2(new_n259), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT7), .A4(G20), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n437), .A2(new_n438), .A3(new_n203), .ZN(new_n439));
  INV_X1    g0239(.A(new_n408), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n436), .B(new_n417), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n253), .A3(new_n413), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n436), .B1(new_n416), .B2(new_n417), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n395), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n430), .A2(new_n323), .A3(new_n431), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n349), .B1(new_n425), .B2(new_n428), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT83), .A3(new_n445), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n435), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n447), .ZN(new_n453));
  INV_X1    g0253(.A(new_n414), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n419), .A2(new_n454), .A3(new_n441), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n453), .A2(KEYINPUT17), .A3(new_n455), .A4(new_n395), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  INV_X1    g0257(.A(new_n433), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n444), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n434), .A2(new_n450), .A3(new_n456), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n337), .A2(G232), .A3(new_n338), .ZN(new_n461));
  INV_X1    g0261(.A(G107), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n461), .B1(new_n462), .B2(new_n337), .C1(new_n341), .C2(new_n215), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n291), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n301), .A2(G244), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n465), .A2(new_n305), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G179), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT74), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT15), .B(G87), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G33), .A3(new_n259), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT73), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n357), .A2(new_n262), .B1(new_n226), .B2(G77), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n472), .A2(KEYINPUT73), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n253), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n272), .A2(G77), .A3(new_n273), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G77), .B2(new_n267), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n467), .A2(new_n388), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n482), .A2(KEYINPUT74), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n469), .B(new_n481), .C1(new_n483), .C2(new_n468), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(G200), .B2(new_n467), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n323), .B2(new_n467), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n392), .A2(new_n460), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT86), .B1(new_n489), .B2(G41), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT86), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n295), .A3(KEYINPUT5), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n207), .B(G45), .C1(new_n295), .C2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n493), .A2(new_n495), .B1(new_n299), .B2(new_n300), .ZN(new_n496));
  OAI211_X1 g0296(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n497));
  OAI211_X1 g0297(.A(G250), .B(new_n338), .C1(new_n283), .C2(new_n284), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n496), .A2(G264), .B1(new_n500), .B2(new_n291), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n304), .A2(new_n493), .A3(new_n495), .A4(G274), .ZN(new_n502));
  AOI21_X1  g0302(.A(G169), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(G179), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n207), .A2(G33), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n370), .A2(new_n371), .A3(new_n267), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n462), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n271), .A2(new_n462), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT25), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT22), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n223), .B(new_n225), .C1(new_n283), .C2(new_n284), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n216), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n462), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n223), .B2(new_n225), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n523), .A2(G20), .B1(new_n520), .B2(new_n462), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n337), .A2(new_n259), .A3(KEYINPUT22), .A4(G87), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT24), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT24), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n519), .A2(new_n525), .A3(new_n529), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n253), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT89), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n516), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n369), .B1(new_n528), .B2(new_n530), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT89), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n506), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n515), .B1(new_n535), .B2(KEYINPUT89), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n500), .A2(new_n291), .ZN(new_n539));
  INV_X1    g0339(.A(new_n493), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(new_n304), .C1(new_n540), .C2(new_n494), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n323), .A2(new_n539), .A3(new_n541), .A4(new_n502), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n349), .B2(new_n505), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n533), .B(new_n369), .C1(new_n528), .C2(new_n530), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n538), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT91), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n501), .A2(new_n502), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n503), .B1(new_n328), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n538), .B2(new_n544), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n532), .A2(new_n533), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n501), .A2(new_n323), .A3(new_n502), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n547), .B2(G200), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n550), .A2(new_n536), .A3(new_n552), .A4(new_n515), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT91), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n546), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n496), .A2(G257), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n502), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G283), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT85), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n337), .A2(new_n563), .A3(G244), .A4(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G244), .B(new_n338), .C1(new_n283), .C2(new_n284), .ZN(new_n567));
  XNOR2_X1  g0367(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n565), .B(G244), .C1(new_n284), .C2(new_n283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT85), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n562), .A2(new_n566), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n291), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n559), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G200), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n437), .A2(new_n438), .A3(new_n462), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n262), .A2(G77), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  INV_X1    g0378(.A(G97), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n578), .A2(new_n579), .A3(G107), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n577), .B1(new_n582), .B2(new_n259), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n253), .B1(new_n576), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n508), .A2(new_n579), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n267), .A2(G97), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n575), .B(new_n589), .C1(new_n323), .C2(new_n574), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n569), .A2(new_n561), .A3(new_n560), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n571), .A2(new_n566), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n290), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n388), .B1(new_n593), .B2(new_n558), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n559), .A2(new_n573), .A3(new_n328), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G264), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n598));
  OAI211_X1 g0398(.A(G257), .B(new_n338), .C1(new_n283), .C2(new_n284), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n337), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n291), .ZN(new_n602));
  OAI211_X1 g0402(.A(G270), .B(new_n304), .C1(new_n540), .C2(new_n494), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n502), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n207), .B2(G33), .ZN(new_n606));
  INV_X1    g0406(.A(G13), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(G1), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n208), .A2(G116), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n272), .A2(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n227), .B2(new_n252), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n257), .A2(G97), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n223), .A2(new_n225), .A3(new_n612), .A4(new_n561), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT20), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n604), .A2(new_n616), .A3(G169), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT88), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(KEYINPUT88), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n616), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n622), .A2(new_n604), .A3(new_n328), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n616), .B1(new_n604), .B2(G200), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n323), .B2(new_n604), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n619), .A2(new_n621), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n223), .A2(new_n225), .A3(G33), .A4(G97), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT19), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n337), .A2(new_n259), .A3(G68), .ZN(new_n631));
  NAND3_X1  g0431(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n223), .A2(new_n225), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n216), .A2(new_n579), .A3(new_n462), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n253), .B1(new_n271), .B2(new_n470), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n508), .A2(new_n216), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(G244), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n640));
  OAI211_X1 g0440(.A(G238), .B(new_n338), .C1(new_n283), .C2(new_n284), .ZN(new_n641));
  NAND2_X1  g0441(.A1(G33), .A2(G116), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n291), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n207), .A2(G45), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n217), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n304), .B(new_n646), .C1(G274), .C2(new_n645), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(G190), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n644), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n639), .A2(new_n650), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n636), .A2(new_n253), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n255), .A2(new_n267), .A3(new_n471), .A4(new_n507), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n470), .A2(new_n271), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n388), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n644), .A2(new_n328), .A3(new_n647), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n597), .A2(new_n627), .A3(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n334), .A2(new_n488), .A3(new_n556), .A4(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n391), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT94), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n420), .B2(new_n433), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n444), .A2(KEYINPUT94), .A3(new_n458), .ZN(new_n668));
  XNOR2_X1  g0468(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n669), .ZN(new_n671));
  AOI211_X1 g0471(.A(new_n666), .B(new_n433), .C1(new_n455), .C2(new_n395), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT94), .B1(new_n444), .B2(new_n458), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n469), .A2(new_n481), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n468), .B1(KEYINPUT74), .B2(new_n482), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n332), .B2(new_n333), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n450), .A2(new_n456), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n281), .A2(new_n317), .A3(new_n324), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n670), .B(new_n674), .C1(new_n678), .C2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n381), .A2(new_n386), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n665), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n488), .A2(new_n334), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n652), .A2(new_n637), .A3(new_n648), .A4(new_n638), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n661), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n596), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT93), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n691), .B(new_n686), .C1(new_n596), .C2(new_n688), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n594), .A2(new_n588), .A3(new_n595), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .A3(new_n661), .A4(new_n654), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n661), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n617), .A2(KEYINPUT88), .A3(new_n620), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n620), .B1(new_n617), .B2(KEYINPUT88), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n697), .A2(new_n698), .A3(new_n623), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT92), .B1(new_n699), .B2(new_n549), .ZN(new_n700));
  INV_X1    g0500(.A(new_n688), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n553), .A2(new_n590), .A3(new_n596), .A4(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n699), .A2(KEYINPUT92), .A3(new_n549), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n684), .B1(new_n685), .B2(new_n708), .ZN(G369));
  NAND2_X1  g0509(.A1(new_n259), .A2(new_n608), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G343), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n534), .B2(new_n536), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n554), .B1(new_n549), .B2(new_n553), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT97), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT97), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n556), .A2(new_n722), .A3(new_n717), .ZN(new_n723));
  INV_X1    g0523(.A(new_n715), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n721), .A2(new_n723), .B1(new_n537), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n619), .A2(new_n621), .A3(new_n624), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n715), .A2(new_n622), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n627), .B2(new_n729), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n727), .B1(new_n731), .B2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n727), .A3(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n537), .A2(new_n715), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n728), .A2(new_n715), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n721), .A2(new_n723), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(G399));
  NAND2_X1  g0541(.A1(new_n211), .A2(new_n295), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n207), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n634), .A2(G116), .ZN(new_n745));
  INV_X1    g0545(.A(new_n231), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n743), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT98), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n661), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n693), .A2(new_n701), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(KEYINPUT26), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n693), .A2(new_n686), .A3(new_n661), .A4(new_n654), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n699), .A2(new_n549), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n753), .B(new_n754), .C1(new_n756), .C2(new_n702), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n749), .B1(new_n757), .B2(new_n715), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n724), .B1(new_n696), .B2(new_n706), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n749), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n556), .A2(new_n663), .A3(new_n715), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT30), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n501), .A2(new_n644), .A3(new_n647), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n604), .A2(new_n328), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n765), .B2(new_n574), .ZN(new_n766));
  INV_X1    g0566(.A(new_n574), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n767), .A2(KEYINPUT30), .A3(new_n764), .A4(new_n763), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n604), .A2(new_n328), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n769), .A2(new_n574), .A3(new_n505), .A4(new_n651), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n724), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT31), .B1(new_n771), .B2(new_n724), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n761), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G330), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n760), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n748), .B1(new_n777), .B2(G1), .ZN(G364));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n731), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n227), .B1(G20), .B2(new_n388), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n323), .A2(new_n349), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G20), .A3(new_n328), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n259), .A2(new_n328), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n323), .A2(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n337), .B1(new_n216), .B2(new_n787), .C1(new_n793), .C2(new_n202), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n226), .A2(new_n328), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G159), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(KEYINPUT32), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n226), .B1(new_n791), .B2(G179), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT103), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G97), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n349), .A2(G190), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n226), .A2(new_n328), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n462), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n788), .A2(new_n808), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n788), .A2(new_n795), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n203), .A2(new_n811), .B1(new_n812), .B2(new_n340), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n788), .A2(new_n786), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n810), .B(new_n813), .C1(G50), .C2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n799), .A2(new_n800), .A3(new_n807), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n399), .B1(new_n787), .B2(new_n600), .C1(new_n809), .C2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G326), .C2(new_n815), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n806), .A2(G294), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n797), .A2(G329), .ZN(new_n824));
  XOR2_X1   g0624(.A(KEYINPUT33), .B(G317), .Z(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT104), .ZN(new_n826));
  INV_X1    g0626(.A(new_n811), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G322), .A2(new_n792), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n785), .B1(new_n817), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n226), .A2(new_n607), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G45), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n744), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n211), .A2(new_n337), .ZN(new_n835));
  INV_X1    g0635(.A(G355), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n835), .A2(new_n836), .B1(G116), .B2(new_n211), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n211), .A2(new_n399), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n296), .B2(new_n746), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT102), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n250), .A2(KEYINPUT101), .A3(new_n296), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT101), .B1(new_n250), .B2(new_n296), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n781), .A2(new_n784), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n834), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n783), .A2(new_n830), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT100), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n735), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n733), .A2(KEYINPUT100), .A3(new_n734), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n731), .A2(G330), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n854), .A2(new_n855), .A3(new_n834), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n848), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT105), .Z(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G396));
  NAND3_X1  g0659(.A1(new_n677), .A2(new_n481), .A3(new_n724), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n724), .A2(new_n481), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n484), .A2(new_n486), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n759), .B(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n834), .B1(new_n864), .B2(new_n776), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n776), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n784), .A2(new_n779), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n834), .B1(G77), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(G294), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n793), .A2(new_n870), .B1(new_n818), .B2(new_n796), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G303), .B2(new_n815), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n399), .B1(new_n787), .B2(new_n462), .ZN(new_n873));
  INV_X1    g0673(.A(new_n812), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(G116), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n809), .A2(new_n216), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n827), .B2(G283), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n872), .A2(new_n807), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n337), .B1(new_n787), .B2(new_n201), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n809), .A2(new_n203), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n879), .B(new_n880), .C1(G132), .C2(new_n797), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT106), .B(G143), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n792), .A2(new_n882), .B1(new_n815), .B2(G137), .ZN(new_n883));
  INV_X1    g0683(.A(G150), .ZN(new_n884));
  INV_X1    g0684(.A(G159), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n883), .B1(new_n884), .B2(new_n811), .C1(new_n885), .C2(new_n812), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT107), .B(KEYINPUT34), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n881), .B1(new_n202), .B2(new_n805), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n869), .B1(new_n890), .B2(new_n784), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n863), .B2(new_n780), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n866), .A2(new_n892), .ZN(G384));
  NOR2_X1   g0693(.A1(new_n831), .A2(new_n207), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n714), .B1(new_n674), .B2(new_n670), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n331), .A2(new_n329), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n330), .B1(new_n316), .B2(G169), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n333), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n333), .A2(new_n724), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n680), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n333), .B(new_n724), .C1(new_n332), .C2(new_n325), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n704), .A2(new_n700), .A3(new_n702), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n695), .A2(new_n661), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n715), .B(new_n863), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n484), .A2(new_n724), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n413), .A2(new_n372), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n399), .A2(new_n259), .A3(new_n400), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(G68), .C1(new_n400), .C2(new_n410), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT16), .B1(new_n912), .B2(new_n408), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n395), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT109), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT109), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n395), .B(new_n916), .C1(new_n910), .C2(new_n913), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n915), .A2(new_n714), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n460), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT37), .B1(new_n444), .B2(new_n458), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n455), .A2(new_n395), .A3(new_n446), .A4(new_n448), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n444), .A2(new_n714), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n429), .ZN(new_n924));
  INV_X1    g0724(.A(new_n432), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(new_n713), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n915), .A2(new_n926), .A3(new_n917), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT37), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n919), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n919), .A2(new_n930), .A3(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n895), .B1(new_n909), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n919), .A2(new_n930), .A3(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n936), .A2(new_n931), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n332), .A2(new_n333), .A3(new_n715), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n674), .A2(new_n679), .A3(new_n670), .ZN(new_n942));
  INV_X1    g0742(.A(new_n922), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n922), .A2(new_n921), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n667), .B2(new_n668), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n923), .B1(new_n946), .B2(new_n929), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT38), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n936), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n939), .B(new_n941), .C1(new_n950), .C2(KEYINPUT39), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n935), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n760), .A2(new_n685), .ZN(new_n953));
  INV_X1    g0753(.A(new_n684), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n952), .B(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(G330), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n775), .A2(new_n902), .A3(new_n863), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT40), .B1(new_n950), .B2(new_n958), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n775), .A2(new_n902), .A3(new_n863), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT40), .B1(new_n932), .B2(new_n933), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n685), .B1(new_n761), .B2(new_n774), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n963), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n894), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n956), .B2(new_n966), .ZN(new_n968));
  INV_X1    g0768(.A(new_n582), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n605), .B(new_n229), .C1(new_n969), .C2(KEYINPUT35), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(KEYINPUT35), .B2(new_n969), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT36), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n746), .A2(G77), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n404), .A2(new_n406), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n973), .A2(new_n974), .B1(G50), .B2(new_n203), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(G1), .A3(new_n607), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT108), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n968), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT110), .ZN(G367));
  NOR2_X1   g0780(.A1(new_n639), .A2(new_n715), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT111), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(new_n661), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n701), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n989));
  INV_X1    g0789(.A(new_n597), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n589), .B2(new_n715), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n693), .A2(new_n724), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n740), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n596), .B1(new_n991), .B2(new_n549), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n715), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n988), .B(new_n989), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n736), .A2(new_n994), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1000), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n995), .A2(KEYINPUT42), .B1(new_n715), .B2(new_n997), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1003), .A2(new_n1004), .A3(new_n987), .A4(new_n986), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n1001), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n742), .B(KEYINPUT41), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n740), .A2(new_n737), .A3(new_n993), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n740), .A2(new_n737), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT44), .B1(new_n1014), .B2(new_n994), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT44), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1016), .B(new_n993), .C1(new_n740), .C2(new_n737), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1012), .A2(new_n1013), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n736), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n537), .A2(new_n724), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n722), .B1(new_n556), .B2(new_n717), .ZN(new_n1022));
  AOI211_X1 g0822(.A(KEYINPUT97), .B(new_n716), .C1(new_n546), .C2(new_n555), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n738), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n740), .B1(new_n1024), .B2(KEYINPUT112), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT112), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n725), .B2(new_n738), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n852), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1024), .A2(KEYINPUT112), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n725), .A2(new_n1026), .A3(new_n738), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1029), .A2(new_n1030), .A3(new_n735), .A4(new_n740), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1028), .A2(new_n777), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n993), .B1(new_n740), .B2(new_n737), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT44), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1010), .B(new_n1011), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n736), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1020), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1009), .B1(new_n1037), .B2(new_n777), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n832), .A2(G1), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1008), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n845), .B1(new_n211), .B2(new_n470), .C1(new_n242), .C2(new_n838), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n834), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n797), .A2(G137), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n793), .B2(new_n884), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G159), .B2(new_n827), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n809), .A2(new_n340), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n787), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n399), .B(new_n1047), .C1(G58), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n806), .A2(G68), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G50), .A2(new_n874), .B1(new_n815), .B2(new_n882), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n787), .A2(new_n605), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT46), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G283), .B2(new_n874), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n870), .A2(new_n811), .B1(new_n814), .B2(new_n818), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G303), .B2(new_n792), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(new_n462), .C2(new_n805), .ZN(new_n1058));
  INV_X1    g0858(.A(G317), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n399), .B1(new_n796), .B2(new_n1059), .C1(new_n579), .C2(new_n809), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT114), .Z(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT47), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n784), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1043), .B1(new_n1065), .B2(new_n1066), .C1(new_n985), .C2(new_n782), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1040), .A2(new_n1067), .ZN(G387));
  NAND3_X1  g0868(.A1(new_n1028), .A2(new_n1039), .A3(new_n1031), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n835), .A2(new_n745), .B1(G107), .B2(new_n211), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n239), .A2(new_n296), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT115), .Z(new_n1072));
  INV_X1    g0872(.A(new_n745), .ZN(new_n1073));
  AOI211_X1 g0873(.A(G45), .B(new_n1073), .C1(G68), .C2(G77), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n356), .A2(G50), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT50), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n838), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1070), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n834), .B1(new_n1078), .B2(new_n846), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n806), .A2(new_n471), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n203), .A2(new_n812), .B1(new_n814), .B2(new_n885), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G150), .B2(new_n797), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n337), .B1(new_n787), .B2(new_n340), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n809), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(G97), .B2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G50), .A2(new_n792), .B1(new_n827), .B2(new_n357), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1080), .A2(new_n1082), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n793), .A2(new_n1059), .B1(new_n600), .B2(new_n812), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT116), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT116), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G311), .A2(new_n827), .B1(new_n815), .B2(G322), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n805), .A2(new_n820), .B1(new_n870), .B2(new_n787), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(KEYINPUT49), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n337), .B1(new_n797), .B2(G326), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n605), .C2(new_n809), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT49), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1087), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1079), .B1(new_n1101), .B2(new_n784), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n726), .B2(new_n782), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1028), .A2(new_n777), .A3(new_n1031), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n743), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n777), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1069), .B(new_n1103), .C1(new_n1105), .C2(new_n1106), .ZN(G393));
  NAND2_X1  g0907(.A1(new_n1020), .A2(new_n1036), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1104), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n743), .A3(new_n1037), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1020), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n247), .A2(new_n211), .A3(new_n399), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n845), .B1(new_n579), .B2(new_n211), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n834), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n870), .A2(new_n812), .B1(new_n811), .B2(new_n600), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G322), .B2(new_n797), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n337), .B(new_n810), .C1(G283), .C2(new_n1048), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n605), .C2(new_n805), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G311), .A2(new_n792), .B1(new_n815), .B2(G317), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT52), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G159), .A2(new_n792), .B1(new_n815), .B2(G150), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT51), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n806), .A2(G77), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n399), .B(new_n876), .C1(G68), .C2(new_n1048), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n827), .A2(G50), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n874), .A2(new_n357), .B1(new_n797), .B2(new_n882), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1118), .A2(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1114), .B1(new_n1128), .B2(new_n784), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n993), .B2(new_n782), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1111), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1110), .A2(new_n1131), .ZN(G390));
  NOR2_X1   g0932(.A1(new_n672), .A2(new_n673), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT37), .B1(new_n1133), .B2(new_n945), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n943), .A2(new_n942), .B1(new_n1134), .B2(new_n923), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n933), .B1(new_n1135), .B2(KEYINPUT38), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n753), .A2(new_n754), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n990), .A2(new_n755), .A3(new_n553), .A4(new_n701), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n724), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n907), .B1(new_n1139), .B2(new_n863), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1136), .B(new_n940), .C1(new_n903), .C2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n938), .B1(new_n1136), .B2(new_n937), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n906), .A2(new_n908), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n941), .B1(new_n1143), .B2(new_n902), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n775), .A2(G330), .A3(new_n863), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(new_n903), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n761), .A2(new_n774), .B1(new_n862), .B2(new_n860), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(G330), .A3(new_n902), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1141), .B(new_n1150), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n775), .A2(new_n488), .A3(G330), .A4(new_n334), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n684), .B(new_n1153), .C1(new_n760), .C2(new_n685), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n902), .B1(new_n1149), .B2(G330), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1143), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1146), .A2(new_n903), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n1150), .A3(new_n1140), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1154), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n742), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1148), .A2(new_n1159), .A3(new_n1151), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1148), .A2(new_n1039), .A3(new_n1151), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n834), .B1(new_n357), .B2(new_n868), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n812), .A2(new_n579), .B1(new_n870), .B2(new_n796), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G283), .B2(new_n815), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n337), .B(new_n880), .C1(G87), .C2(new_n1048), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G116), .A2(new_n792), .B1(new_n827), .B2(G107), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1123), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G132), .A2(new_n792), .B1(new_n815), .B2(G128), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT117), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n806), .A2(G159), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n399), .B1(new_n1084), .B2(G50), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT54), .B(G143), .Z(new_n1176));
  NAND3_X1  g0976(.A1(new_n1048), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT53), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n787), .B2(new_n884), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n874), .A2(new_n1176), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n827), .A2(G137), .B1(G125), .B2(new_n797), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1174), .A2(new_n1175), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1171), .B1(new_n1173), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1166), .B1(new_n1183), .B2(new_n784), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1142), .B2(new_n780), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1164), .A2(new_n1165), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1165), .B1(new_n1164), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1163), .B1(new_n1186), .B2(new_n1187), .ZN(G378));
  NAND2_X1  g0988(.A1(new_n935), .A2(new_n951), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n382), .A2(new_n714), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n392), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n381), .A2(new_n386), .A3(new_n391), .A4(new_n1190), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1195), .A2(new_n1196), .A3(KEYINPUT121), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n963), .B2(G330), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n957), .B(new_n1197), .C1(new_n959), .C2(new_n962), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1189), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT38), .B1(new_n944), .B2(new_n947), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n902), .B(new_n1149), .C1(new_n1202), .C2(new_n936), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1203), .A2(KEYINPUT40), .B1(new_n960), .B2(new_n961), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1197), .B1(new_n1204), .B2(new_n957), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n963), .A2(G330), .A3(new_n1198), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n952), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1039), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n792), .A2(G107), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1050), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n337), .A2(G41), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n340), .B2(new_n787), .C1(new_n814), .C2(new_n605), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G58), .A2(new_n1084), .B1(new_n797), .B2(G283), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n579), .B2(new_n811), .C1(new_n470), .C2(new_n812), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1219), .C1(new_n1213), .C2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n257), .B(new_n295), .C1(new_n809), .C2(new_n885), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n874), .A2(G137), .B1(new_n1048), .B2(new_n1176), .ZN(new_n1223));
  INV_X1    g1023(.A(G128), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n793), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G132), .B2(new_n827), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n806), .A2(G150), .B1(G125), .B2(new_n815), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT120), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1223), .B(new_n1226), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1222), .B(new_n1232), .C1(G124), .C2(new_n797), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1221), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n834), .B1(G50), .B2(new_n868), .C1(new_n1235), .C2(new_n785), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1195), .A2(new_n1196), .A3(new_n780), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1209), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1154), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1201), .A2(new_n1207), .B1(new_n1162), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n742), .B1(new_n1242), .B2(KEYINPUT57), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1162), .A2(new_n1241), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1208), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT57), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1240), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(G375));
  AOI22_X1  g1049(.A1(new_n1156), .A2(new_n1158), .B1(G1), .B2(new_n832), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT122), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT122), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n834), .B1(G68), .B2(new_n868), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n462), .A2(new_n812), .B1(new_n814), .B2(new_n870), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G303), .B2(new_n797), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n337), .B(new_n1047), .C1(G97), .C2(new_n1048), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G283), .A2(new_n792), .B1(new_n827), .B2(G116), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1080), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n806), .A2(G50), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n399), .B1(new_n1084), .B2(G58), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G137), .A2(new_n792), .B1(new_n827), .B2(new_n1176), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G132), .A2(new_n815), .B1(new_n874), .B2(G150), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n796), .A2(new_n1224), .B1(new_n885), .B2(new_n787), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT123), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1258), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1253), .B1(new_n1266), .B2(new_n784), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n902), .B2(new_n780), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1251), .A2(new_n1252), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1009), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1156), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1160), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(G381));
  NAND2_X1  g1073(.A1(new_n1164), .A2(new_n1185), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1277), .A2(G390), .A3(G381), .A4(G384), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1278), .A2(new_n1040), .A3(new_n1067), .A4(new_n1248), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT124), .Z(G407));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1275), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(G343), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1248), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G407), .A2(new_n1284), .ZN(G409));
  AOI21_X1  g1085(.A(new_n1238), .B1(new_n1208), .B2(new_n1039), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1208), .A2(KEYINPUT57), .A3(new_n1244), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n743), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1242), .A2(KEYINPUT57), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1286), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1245), .A2(new_n1009), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1275), .B1(new_n1291), .B2(new_n1240), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1281), .A2(G343), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1271), .B1(new_n1159), .B2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1156), .A2(new_n1154), .A3(KEYINPUT60), .A4(new_n1158), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n743), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1269), .A2(G384), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1297), .A2(new_n743), .A3(new_n1298), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1251), .A2(new_n1252), .A3(new_n1268), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1293), .A2(new_n1295), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1294), .A2(G2897), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1305), .B(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1293), .A2(new_n1313), .A3(new_n1295), .A4(new_n1306), .ZN(new_n1314));
  XOR2_X1   g1114(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1315));
  NAND4_X1  g1115(.A1(new_n1308), .A2(new_n1312), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1040), .A2(G390), .A3(new_n1067), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT126), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(G393), .B(new_n858), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(G390), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G387), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1317), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1322), .A2(new_n1319), .A3(new_n1325), .A4(new_n1317), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1316), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1326), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1318), .A2(new_n1319), .B1(new_n1322), .B2(new_n1317), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1329), .A2(new_n1330), .A3(KEYINPUT61), .ZN(new_n1331));
  AOI211_X1 g1131(.A(new_n1294), .B(new_n1305), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT125), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT63), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1307), .A2(KEYINPUT125), .A3(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1331), .A2(new_n1312), .A3(new_n1334), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1328), .A2(new_n1337), .ZN(G405));
  OAI21_X1  g1138(.A(new_n1290), .B1(new_n1248), .B2(new_n1282), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1329), .A2(new_n1330), .A3(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1339), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1305), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1327), .A2(new_n1340), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1324), .A2(new_n1326), .A3(new_n1339), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(new_n1306), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1343), .A2(new_n1346), .ZN(G402));
endmodule


