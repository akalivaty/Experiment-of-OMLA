//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT94), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(new_n203), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT21), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT95), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G183gat), .B(G211gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(KEYINPUT16), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n217), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT89), .B(G8gat), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n222), .A2(KEYINPUT90), .B1(new_n223), .B2(new_n220), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n222), .A2(KEYINPUT90), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT91), .B1(new_n224), .B2(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231));
  INV_X1    g030(.A(new_n210), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G127gat), .B(G155gat), .Z(new_n234));
  NAND2_X1  g033(.A1(G231gat), .A2(G233gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n233), .A2(new_n236), .ZN(new_n238));
  OR3_X1    g037(.A1(new_n216), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n216), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G43gat), .B(G50gat), .Z(new_n242));
  INV_X1    g041(.A(G29gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n244));
  INV_X1    g043(.A(G36gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n243), .B2(KEYINPUT14), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT14), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G29gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n242), .B1(new_n249), .B2(KEYINPUT15), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(KEYINPUT15), .B2(new_n249), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(KEYINPUT15), .A3(new_n242), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT7), .ZN(new_n256));
  NAND2_X1  g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257));
  INV_X1    g056(.A(G85gat), .ZN(new_n258));
  INV_X1    g057(.A(G92gat), .ZN(new_n259));
  AOI22_X1  g058(.A1(KEYINPUT8), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G99gat), .B(G106gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT97), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT98), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n254), .A2(KEYINPUT98), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G232gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n253), .A2(new_n263), .B1(KEYINPUT41), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n273), .A3(new_n275), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n272), .A2(KEYINPUT41), .ZN(new_n279));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n281), .B(KEYINPUT96), .Z(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT99), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n278), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n275), .B1(new_n270), .B2(new_n273), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n281), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n283), .A3(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT100), .B1(new_n263), .B2(new_n210), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n210), .B2(new_n263), .ZN(new_n293));
  INV_X1    g092(.A(new_n263), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n232), .A3(KEYINPUT100), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT10), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT10), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n294), .A2(new_n232), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n291), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(new_n295), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G176gat), .B(G204gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n241), .A2(new_n290), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT93), .ZN(new_n311));
  XOR2_X1   g110(.A(G15gat), .B(G43gat), .Z(new_n312));
  XNOR2_X1  g111(.A(G71gat), .B(G99gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G183gat), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT28), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(KEYINPUT26), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n330), .A2(new_n331), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n323), .A2(new_n317), .A3(new_n319), .A4(new_n320), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n325), .A2(new_n329), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT64), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n338), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT64), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(G169gat), .B2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n327), .A2(KEYINPUT65), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT65), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G169gat), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT23), .A4(new_n328), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n342), .A2(new_n343), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n334), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  NAND2_X1  g157(.A1(G113gat), .A2(G120gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G127gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G134gat), .ZN(new_n362));
  INV_X1    g161(.A(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G127gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n354), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT1), .B1(new_n355), .B2(new_n356), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n367), .A2(KEYINPUT70), .A3(new_n359), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT69), .B1(new_n363), .B2(G127gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT69), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n361), .A3(G134gat), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT68), .B(G134gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G127gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n371), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n336), .A2(new_n335), .B1(new_n380), .B2(G190gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT23), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n345), .A3(new_n346), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT25), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n353), .A2(KEYINPUT71), .A3(new_n379), .A4(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT71), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n334), .A2(new_n352), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT68), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G134gat), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n388), .A2(new_n390), .A3(G127gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n374), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n360), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n366), .A3(new_n369), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n386), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n387), .A2(new_n394), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n385), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n315), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n397), .B2(new_n399), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI221_X4 g205(.A(new_n403), .B1(KEYINPUT33), .B2(new_n314), .C1(new_n397), .C2(new_n399), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT34), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n398), .B2(KEYINPUT73), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n385), .A2(new_n398), .A3(new_n395), .A4(new_n396), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n413), .A2(KEYINPUT74), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(KEYINPUT74), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n387), .A2(new_n394), .A3(new_n386), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n387), .A2(new_n394), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT74), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n398), .A4(new_n395), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n413), .A2(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n411), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT76), .B1(new_n409), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n421), .A2(new_n411), .A3(new_n422), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n411), .B1(new_n421), .B2(new_n422), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT76), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n408), .A4(new_n406), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT36), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n409), .A2(new_n424), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT33), .B1(new_n397), .B2(new_n399), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n404), .A2(new_n435), .A3(new_n315), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT72), .B1(new_n436), .B2(new_n407), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n406), .A2(new_n408), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n439), .A3(new_n424), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT75), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT75), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .A4(new_n424), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n431), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n434), .B1(KEYINPUT36), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G197gat), .B(G204gat), .ZN(new_n446));
  INV_X1    g245(.A(G211gat), .ZN(new_n447));
  INV_X1    g246(.A(G218gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(KEYINPUT22), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G211gat), .B(G218gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n387), .A2(G226gat), .A3(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT29), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n387), .A2(new_n454), .B1(G226gat), .B2(G233gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n387), .A2(new_n454), .ZN(new_n457));
  NAND2_X1  g256(.A1(G226gat), .A2(G233gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n452), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n387), .A2(G226gat), .A3(G233gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  NAND4_X1  g264(.A1(new_n456), .A2(new_n462), .A3(KEYINPUT30), .A4(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT77), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n456), .B2(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n462), .A3(new_n465), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n475), .B2(KEYINPUT2), .ZN(new_n476));
  XNOR2_X1  g275(.A(G141gat), .B(G148gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT2), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(new_n474), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT80), .B1(new_n483), .B2(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n481), .A2(new_n474), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT2), .B1(new_n477), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT79), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n487), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n379), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n394), .B1(new_n493), .B2(new_n485), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT81), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OR3_X1    g300(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n477), .A2(new_n488), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n482), .A3(new_n492), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n486), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n484), .A4(new_n480), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT3), .B1(new_n485), .B2(new_n493), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n394), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n484), .A3(new_n480), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n394), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n494), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n509), .A2(new_n512), .A3(new_n501), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n498), .A2(KEYINPUT82), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n502), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G1gat), .B(G29gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT0), .ZN(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G85gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524));
  INV_X1    g323(.A(new_n522), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n502), .C1(new_n516), .C2(new_n517), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n518), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n525), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n472), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n460), .B1(new_n507), .B2(new_n454), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n506), .B1(new_n452), .B2(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n511), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  NAND2_X1  g334(.A1(G228gat), .A2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G22gat), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G50gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n535), .B(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n530), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT83), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n495), .A2(new_n542), .A3(new_n501), .A4(new_n496), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n543), .A2(KEYINPUT39), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n500), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n495), .A2(new_n501), .A3(new_n496), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT83), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT39), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n550), .A3(new_n500), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n549), .A2(KEYINPUT40), .A3(new_n522), .A4(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n552), .A2(new_n526), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT40), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n522), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT84), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT84), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n553), .A2(new_n558), .A3(new_n472), .A4(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(new_n540), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n527), .A2(new_n529), .ZN(new_n563));
  INV_X1    g362(.A(new_n469), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n456), .A2(new_n462), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT85), .B1(new_n565), .B2(KEYINPUT37), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT85), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n456), .A2(new_n462), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n465), .B1(new_n565), .B2(KEYINPUT37), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n564), .B1(new_n572), .B2(KEYINPUT38), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT86), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT86), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n577), .A3(new_n574), .A4(new_n571), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n563), .A2(new_n573), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n541), .B1(new_n562), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n441), .A2(new_n431), .A3(new_n540), .A4(new_n443), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n527), .A2(new_n529), .ZN(new_n582));
  INV_X1    g381(.A(new_n472), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT35), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n425), .A2(new_n430), .B1(new_n409), .B2(new_n424), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n530), .A3(new_n587), .A4(new_n540), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n445), .A2(new_n580), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n228), .A2(new_n229), .A3(new_n253), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n254), .A2(new_n226), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n591), .ZN(new_n598));
  INV_X1    g397(.A(new_n590), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n253), .B1(new_n228), .B2(new_n229), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT88), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G113gat), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G141gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n601), .A4(new_n609), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n311), .B1(new_n589), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n585), .A2(new_n588), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n572), .A2(KEYINPUT38), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n527), .A2(new_n618), .A3(new_n529), .A4(new_n469), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n576), .A2(new_n578), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n540), .B(new_n561), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n586), .A2(new_n432), .ZN(new_n622));
  INV_X1    g421(.A(new_n540), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n584), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n617), .A2(new_n621), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(KEYINPUT93), .A3(new_n613), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n310), .B1(new_n615), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n563), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  INV_X1    g429(.A(new_n628), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n631), .A2(new_n583), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n223), .B1(new_n628), .B2(new_n472), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(KEYINPUT42), .B2(new_n633), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n631), .B2(new_n445), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n431), .A2(new_n433), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n638), .A2(G15gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n631), .B2(new_n639), .ZN(G1326gat));
  NAND2_X1  g439(.A1(new_n628), .A2(new_n623), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT101), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(KEYINPUT101), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT43), .B(G22gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(G1327gat));
  AND2_X1   g448(.A1(new_n239), .A2(new_n240), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n285), .A2(new_n289), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n309), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT102), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n615), .A2(new_n627), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n243), .A4(new_n563), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AND4_X1   g457(.A1(new_n617), .A2(new_n622), .A3(new_n621), .A4(new_n624), .ZN(new_n659));
  AOI22_X1  g458(.A1(KEYINPUT75), .A2(new_n440), .B1(new_n425), .B2(new_n430), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n660), .A2(new_n530), .A3(new_n540), .A4(new_n443), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n638), .A2(new_n623), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n661), .A2(KEYINPUT35), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT105), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n616), .A2(new_n666), .A3(new_n625), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n290), .A2(KEYINPUT44), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT106), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n290), .B1(new_n616), .B2(new_n625), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n674), .B(KEYINPUT44), .C1(new_n589), .C2(new_n290), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n665), .A2(new_n677), .A3(new_n667), .A4(new_n668), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n670), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n241), .A2(new_n614), .A3(new_n308), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(new_n563), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n658), .B1(new_n243), .B2(new_n681), .ZN(G1328gat));
  NAND4_X1  g481(.A1(new_n654), .A2(new_n655), .A3(new_n245), .A4(new_n472), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT46), .Z(new_n684));
  NAND3_X1  g483(.A1(new_n679), .A2(new_n472), .A3(new_n680), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G36gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691));
  INV_X1    g490(.A(new_n445), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n679), .A2(new_n692), .A3(new_n680), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n638), .A2(G43gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n654), .A2(new_n655), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n691), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n696), .ZN(new_n698));
  AOI211_X1 g497(.A(KEYINPUT47), .B(new_n698), .C1(new_n693), .C2(G43gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n679), .A2(G50gat), .A3(new_n623), .A4(new_n680), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n654), .A2(new_n623), .A3(new_n655), .ZN(new_n702));
  INV_X1    g501(.A(G50gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT48), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n707), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1331gat));
  AND2_X1   g508(.A1(new_n665), .A2(new_n667), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n650), .A2(new_n651), .A3(new_n613), .A4(new_n309), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n563), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g514(.A1(new_n583), .A2(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n583), .A2(KEYINPUT108), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  AND2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(G1333gat));
  XNOR2_X1  g523(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n586), .A3(new_n711), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n205), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n445), .A2(new_n205), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n711), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT109), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n730), .A2(KEYINPUT109), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n726), .B(new_n728), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n731), .ZN(new_n734));
  INV_X1    g533(.A(new_n728), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n725), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n733), .A2(new_n736), .ZN(G1334gat));
  NOR2_X1   g536(.A1(new_n712), .A2(new_n540), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n206), .ZN(G1335gat));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n671), .A2(new_n614), .A3(new_n650), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n650), .A2(new_n614), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n589), .A2(new_n290), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n743), .A2(new_n746), .B1(new_n742), .B2(new_n741), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(new_n258), .A3(new_n563), .A4(new_n308), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n744), .A2(new_n309), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n679), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(new_n563), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n752), .B2(new_n258), .ZN(G1336gat));
  NAND3_X1  g552(.A1(new_n679), .A2(new_n718), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n718), .A2(new_n259), .A3(new_n308), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT112), .Z(new_n757));
  NAND2_X1  g556(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n746), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n745), .B2(KEYINPUT51), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n741), .A2(KEYINPUT114), .A3(new_n742), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n757), .B(KEYINPUT113), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n760), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n679), .A2(new_n472), .A3(new_n750), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n759), .A2(new_n760), .B1(new_n767), .B2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(G99gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n771), .A3(new_n586), .A4(new_n308), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n751), .A2(new_n692), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n771), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n679), .A2(new_n623), .A3(new_n750), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n309), .A2(G106gat), .A3(new_n540), .ZN(new_n776));
  AOI22_X1  g575(.A1(G106gat), .A2(new_n775), .B1(new_n765), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n775), .A2(G106gat), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n780));
  INV_X1    g579(.A(new_n776), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n747), .B2(new_n781), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n777), .A2(new_n778), .B1(new_n779), .B2(new_n782), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n310), .A2(new_n613), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n305), .B1(new_n299), .B2(KEYINPUT54), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n298), .B1(new_n300), .B2(new_n297), .ZN(new_n788));
  INV_X1    g587(.A(new_n291), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(KEYINPUT54), .A3(new_n299), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n785), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n787), .C2(new_n791), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n791), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n306), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n599), .A2(new_n600), .A3(new_n598), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n608), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n612), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(new_n651), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n794), .ZN(new_n805));
  INV_X1    g604(.A(new_n797), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n792), .A2(new_n785), .A3(new_n793), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n285), .A2(new_n289), .A3(new_n803), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n803), .A2(new_n308), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n798), .B2(new_n613), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n804), .B(new_n810), .C1(new_n813), .C2(new_n651), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n784), .B1(new_n814), .B2(new_n650), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n718), .A2(new_n582), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n581), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n613), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n818), .A2(new_n662), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n614), .A2(new_n355), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G1340gat));
  AOI21_X1  g624(.A(G120gat), .B1(new_n821), .B2(new_n308), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n309), .A2(new_n356), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n823), .B2(new_n827), .ZN(G1341gat));
  AND3_X1   g627(.A1(new_n818), .A2(new_n662), .A3(new_n241), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n241), .A2(new_n361), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n829), .A2(new_n361), .B1(new_n820), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI221_X1 g632(.A(KEYINPUT118), .B1(new_n820), .B2(new_n830), .C1(new_n829), .C2(new_n361), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1342gat));
  NAND2_X1  g634(.A1(new_n814), .A2(new_n650), .ZN(new_n836));
  INV_X1    g635(.A(new_n784), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n582), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n290), .A2(new_n472), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n376), .A3(new_n819), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT56), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n823), .A2(new_n651), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n363), .B2(new_n844), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n836), .A2(new_n837), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n623), .ZN(new_n848));
  XNOR2_X1  g647(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n790), .A2(KEYINPUT54), .A3(new_n299), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n786), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n796), .A4(new_n306), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n613), .ZN(new_n854));
  INV_X1    g653(.A(new_n849), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n787), .B2(new_n791), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT120), .B1(new_n797), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n812), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n810), .B(new_n804), .C1(new_n858), .C2(new_n651), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n784), .B1(new_n859), .B2(new_n650), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n860), .B2(new_n540), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n692), .A2(new_n817), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n848), .A2(new_n861), .A3(new_n613), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G141gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n614), .A2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n445), .A2(new_n623), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n838), .B2(new_n868), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n815), .A2(KEYINPUT121), .A3(new_n582), .A4(new_n867), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n719), .B(new_n865), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n839), .A2(new_n867), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n614), .A2(new_n718), .A3(G141gat), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n863), .A2(G141gat), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n872), .B2(new_n876), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n309), .A2(G148gat), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n719), .B(new_n878), .C1(new_n869), .C2(new_n870), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n848), .A2(new_n861), .A3(new_n862), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n309), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G148gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n540), .A2(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n857), .A2(new_n613), .A3(new_n853), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n651), .B1(new_n886), .B2(new_n811), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n808), .A2(new_n809), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n798), .A2(new_n651), .A3(new_n803), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n890), .B(new_n891), .C1(new_n858), .C2(new_n651), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n889), .A2(new_n892), .A3(new_n650), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n885), .B1(new_n893), .B2(new_n784), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n815), .B2(new_n540), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n894), .A2(new_n308), .A3(new_n862), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n882), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n879), .B1(new_n884), .B2(new_n897), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n241), .A2(G155gat), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT123), .Z(new_n900));
  NOR2_X1   g699(.A1(new_n880), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(G155gat), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n241), .B(new_n719), .C1(new_n869), .C2(new_n870), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n880), .B2(new_n290), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n869), .A2(new_n870), .ZN(new_n906));
  INV_X1    g705(.A(G162gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n840), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n563), .A2(new_n583), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n662), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n815), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n614), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n815), .A2(new_n563), .A3(new_n719), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n819), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n613), .A2(new_n348), .A3(new_n350), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1348gat));
  OAI21_X1  g716(.A(G176gat), .B1(new_n912), .B2(new_n309), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n308), .A2(new_n328), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n915), .B2(new_n919), .ZN(G1349gat));
  NOR3_X1   g719(.A1(new_n815), .A2(new_n650), .A3(new_n911), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n922));
  OAI21_X1  g721(.A(G183gat), .B1(new_n921), .B2(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n241), .A2(new_n317), .A3(new_n319), .ZN(new_n924));
  OAI22_X1  g723(.A1(new_n922), .A2(new_n923), .B1(new_n915), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT60), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  OAI221_X1 g726(.A(new_n927), .B1(new_n915), .B2(new_n924), .C1(new_n922), .C2(new_n923), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1350gat));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  INV_X1    g729(.A(new_n915), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n290), .A2(G190gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR4_X1   g732(.A1(new_n915), .A2(KEYINPUT125), .A3(G190gat), .A4(new_n290), .ZN(new_n934));
  OAI21_X1  g733(.A(G190gat), .B1(new_n912), .B2(new_n290), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n937));
  OAI22_X1  g736(.A1(new_n933), .A2(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  AND2_X1   g737(.A1(new_n914), .A2(new_n868), .ZN(new_n939));
  AOI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n613), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n894), .A2(new_n895), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n445), .A2(new_n910), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n613), .A2(G197gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  NAND3_X1  g745(.A1(new_n941), .A2(new_n308), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G204gat), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  AOI211_X1 g748(.A(G204gat), .B(new_n309), .C1(new_n949), .C2(KEYINPUT62), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n914), .A2(new_n868), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n447), .A3(new_n241), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n894), .A2(new_n241), .A3(new_n895), .A4(new_n943), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n651), .A3(new_n943), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G218gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n448), .A3(new_n651), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


