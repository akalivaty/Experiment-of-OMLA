//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND2_X1  g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AND2_X1   g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(KEYINPUT66), .B1(G567), .B2(new_n456), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n460), .B1(KEYINPUT66), .B2(new_n459), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n467), .A2(G136), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  MUX2_X1   g058(.A(G100), .B(G112), .S(G2105), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OR2_X1    g062(.A1(new_n464), .A2(new_n465), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n488), .A2(G126), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n490), .B2(new_n468), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(KEYINPUT4), .B(G138), .C1(new_n464), .C2(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(G102), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(new_n468), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n488), .A2(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n495), .A2(new_n481), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n501), .A3(KEYINPUT5), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(new_n506), .ZN(new_n521));
  INV_X1    g096(.A(new_n502), .ZN(new_n522));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI211_X1 g102(.A(G51), .B(G543), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n531), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  AND4_X1   g109(.A1(G89), .A2(new_n521), .A3(new_n522), .A4(new_n515), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n520), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(G89), .A3(new_n515), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n533), .A2(new_n528), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT71), .A4(new_n525), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n507), .A2(new_n515), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  INV_X1    g118(.A(new_n513), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT72), .B1(new_n546), .B2(new_n509), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n521), .A2(G64), .A3(new_n522), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(new_n551), .A3(G651), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n545), .B1(new_n547), .B2(new_n552), .ZN(G171));
  NAND3_X1  g128(.A1(new_n521), .A2(G56), .A3(new_n522), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n509), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n521), .A2(G81), .A3(new_n522), .A4(new_n515), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n513), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  XOR2_X1   g138(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n565), .B(new_n566), .Z(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G188));
  NAND3_X1  g143(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n513), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n507), .A2(G91), .A3(new_n515), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n573), .B(new_n574), .C1(new_n509), .C2(new_n575), .ZN(G299));
  INV_X1    g151(.A(new_n545), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n551), .B1(new_n550), .B2(G651), .ZN(new_n578));
  AOI211_X1 g153(.A(KEYINPUT72), .B(new_n509), .C1(new_n548), .C2(new_n549), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n513), .A2(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n516), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n521), .A2(new_n522), .ZN(new_n586));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n509), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n507), .A2(KEYINPUT76), .A3(G61), .ZN(new_n591));
  INV_X1    g166(.A(G73), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n501), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT76), .B1(new_n507), .B2(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n516), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G86), .B1(G48), .B2(new_n513), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n509), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n507), .A2(G85), .A3(new_n515), .ZN(new_n601));
  XOR2_X1   g176(.A(KEYINPUT77), .B(G47), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n513), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT78), .B1(new_n601), .B2(new_n603), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(G290));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(G301), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n507), .A2(G92), .A3(new_n515), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT79), .B(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n586), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(KEYINPUT80), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(KEYINPUT80), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n610), .B1(new_n621), .B2(new_n609), .ZN(G321));
  XNOR2_X1  g197(.A(G321), .B(KEYINPUT81), .ZN(G284));
  NAND2_X1  g198(.A1(G299), .A2(new_n609), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n621), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(new_n560), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n619), .A2(new_n627), .A3(new_n620), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G323));
  XOR2_X1   g207(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n633));
  XNOR2_X1  g208(.A(G323), .B(new_n633), .ZN(G282));
  NAND2_X1  g209(.A1(new_n467), .A2(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  MUX2_X1   g215(.A(G99), .B(G111), .S(G2105), .Z(new_n641));
  AOI22_X1  g216(.A1(new_n482), .A2(G123), .B1(G2104), .B2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  INV_X1    g218(.A(new_n467), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G2096), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n640), .A3(new_n647), .ZN(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2427), .ZN(new_n652));
  INV_X1    g227(.A(G2430), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(G401));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(KEYINPUT85), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(KEYINPUT85), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n668), .B(KEYINPUT17), .Z(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n673), .C1(new_n674), .C2(new_n667), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n667), .A3(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n666), .A3(new_n668), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n646), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2100), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n689), .B1(new_n684), .B2(new_n687), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n692), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  INV_X1    g277(.A(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT91), .B1(new_n703), .B2(G16), .ZN(new_n704));
  OR3_X1    g279(.A1(new_n703), .A2(KEYINPUT91), .A3(G16), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(G166), .C2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(G23), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n589), .B2(new_n706), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n595), .A2(new_n597), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G6), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n702), .B(new_n713), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n706), .A2(G24), .ZN(new_n726));
  XOR2_X1   g301(.A(G290), .B(KEYINPUT89), .Z(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G25), .A2(G29), .ZN(new_n731));
  MUX2_X1   g306(.A(G95), .B(G107), .S(G2105), .Z(new_n732));
  AOI22_X1  g307(.A1(new_n482), .A2(G119), .B1(G2104), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G131), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n644), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n731), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n730), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n725), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n716), .B(new_n717), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(new_n720), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(new_n722), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n702), .B1(new_n748), .B2(new_n713), .ZN(new_n749));
  OAI21_X1  g324(.A(KEYINPUT36), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n713), .B1(new_n723), .B2(new_n724), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT34), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n752), .A2(new_n753), .A3(new_n725), .A4(new_n744), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n467), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n482), .A2(G129), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n469), .A2(G105), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT26), .Z(new_n760));
  NAND4_X1  g335(.A1(new_n756), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n763), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT97), .ZN(new_n768));
  NAND2_X1  g343(.A1(G160), .A2(G29), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n763), .B1(new_n770), .B2(G34), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n771), .A2(KEYINPUT95), .B1(new_n770), .B2(G34), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT95), .B2(new_n771), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT96), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(G2084), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n765), .A2(new_n766), .ZN(new_n777));
  AND2_X1   g352(.A1(KEYINPUT30), .A2(G28), .ZN(new_n778));
  NOR2_X1   g353(.A1(KEYINPUT30), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n763), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n780), .B(new_n782), .C1(new_n645), .C2(new_n763), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n763), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n467), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n482), .A2(G128), .ZN(new_n788));
  MUX2_X1   g363(.A(G104), .B(G116), .S(G2105), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2104), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2067), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n763), .A2(G35), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT100), .Z(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n763), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n784), .B(new_n793), .C1(new_n798), .C2(G2090), .ZN(new_n799));
  AOI21_X1  g374(.A(G2084), .B1(new_n769), .B2(new_n774), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n763), .A2(G27), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n499), .B2(G29), .ZN(new_n803));
  INV_X1    g378(.A(G2078), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n776), .A2(new_n799), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n706), .A2(G4), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n621), .B2(new_n706), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1348), .Z(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G19), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n560), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n469), .A2(G103), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n467), .A2(G139), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n815), .B(new_n816), .C1(new_n481), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT94), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G29), .ZN(new_n820));
  NOR2_X1   g395(.A1(G29), .A2(G33), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT92), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2072), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G21), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G168), .B2(G16), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G1966), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(G1966), .ZN(new_n828));
  AND4_X1   g403(.A1(new_n812), .A2(new_n824), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n798), .A2(KEYINPUT102), .A3(G2090), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT102), .B1(new_n798), .B2(G2090), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n706), .A2(G5), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G171), .B2(new_n706), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G1961), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n706), .A2(G20), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT23), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n573), .A2(new_n574), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n575), .A2(new_n509), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n837), .B1(new_n840), .B2(new_n706), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1956), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n831), .A2(new_n832), .A3(new_n835), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n806), .A2(new_n809), .A3(new_n829), .A4(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT103), .B1(new_n755), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n847));
  AOI211_X1 g422(.A(new_n847), .B(new_n844), .C1(new_n750), .C2(new_n754), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n755), .A2(new_n845), .ZN(G150));
  NAND2_X1  g425(.A1(new_n621), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT105), .B1(new_n556), .B2(new_n559), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n521), .A2(G67), .A3(new_n522), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n509), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n521), .A2(G93), .A3(new_n522), .A4(new_n515), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n513), .A2(G55), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n856), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n507), .B2(G67), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n859), .B(new_n858), .C1(new_n864), .C2(new_n509), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n560), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n862), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n853), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  NAND2_X1  g450(.A1(new_n819), .A2(KEYINPUT106), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n761), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n467), .A2(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n482), .A2(G130), .ZN(new_n880));
  MUX2_X1   g455(.A(G106), .B(G118), .S(G2105), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G2104), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n737), .A2(new_n738), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n636), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n636), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n884), .A2(new_n636), .ZN(new_n889));
  INV_X1    g464(.A(new_n883), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(new_n791), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n499), .B(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n888), .B2(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n878), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n877), .A3(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G160), .B(new_n486), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n645), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n897), .A2(new_n901), .A3(new_n904), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n618), .A2(new_n840), .ZN(new_n911));
  NAND3_X1  g486(.A1(G299), .A2(new_n613), .A3(new_n617), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  NAND4_X1  g492(.A1(G299), .A2(new_n613), .A3(new_n617), .A4(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n911), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n867), .A2(new_n854), .ZN(new_n921));
  INV_X1    g496(.A(new_n862), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n631), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n631), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G305), .A2(G303), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n595), .A2(G166), .A3(new_n597), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G290), .A2(G288), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n589), .B(new_n600), .C1(new_n606), .C2(new_n607), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n631), .A2(new_n923), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n916), .A2(new_n911), .A3(new_n918), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n924), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n927), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n927), .B2(new_n944), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n946), .A2(new_n947), .B1(new_n937), .B2(new_n938), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n942), .A2(new_n943), .A3(new_n924), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n942), .A2(new_n924), .B1(new_n915), .B2(new_n919), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n940), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n937), .A2(new_n938), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n945), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n609), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n865), .A2(G868), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(G295));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  OR3_X1    g532(.A1(new_n954), .A2(new_n957), .A3(new_n955), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G331));
  INV_X1    g535(.A(new_n936), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n536), .B2(new_n539), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G171), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n536), .A2(new_n962), .A3(new_n539), .ZN(new_n965));
  NAND2_X1  g540(.A1(G301), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n923), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n523), .B(new_n502), .C1(new_n504), .C2(new_n506), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n533), .A2(new_n528), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT71), .B1(new_n971), .B2(new_n537), .ZN(new_n972));
  AND4_X1   g547(.A1(KEYINPUT71), .A2(new_n537), .A3(new_n538), .A4(new_n525), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT110), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(G301), .A3(new_n965), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n868), .A2(new_n975), .A3(new_n964), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n968), .A2(new_n976), .B1(new_n915), .B2(new_n919), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n968), .A2(new_n943), .A3(new_n976), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n968), .A2(new_n980), .A3(new_n943), .A4(new_n976), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n961), .B(new_n977), .C1(new_n979), .C2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n868), .A2(new_n975), .A3(new_n964), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n975), .A2(new_n964), .B1(new_n921), .B2(new_n922), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT41), .B(new_n913), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n961), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n968), .A2(new_n976), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n943), .B1(new_n987), .B2(KEYINPUT41), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n907), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n979), .A2(new_n981), .ZN(new_n993));
  INV_X1    g568(.A(new_n977), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n961), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n936), .A3(new_n994), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n907), .A4(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n982), .C2(new_n989), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n992), .A2(KEYINPUT44), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(KEYINPUT43), .A3(new_n907), .A4(new_n998), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n982), .B2(new_n989), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(KEYINPUT113), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(G397));
  NAND4_X1  g585(.A1(new_n478), .A2(G40), .A3(new_n470), .A4(new_n474), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n475), .A2(KEYINPUT114), .A3(G40), .A4(new_n478), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n492), .B2(new_n498), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(KEYINPUT45), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n884), .A2(new_n742), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n884), .A2(new_n742), .ZN(new_n1022));
  INV_X1    g597(.A(G1996), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n761), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2067), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n791), .B(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1022), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G290), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n729), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n729), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT115), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1019), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1017), .A2(KEYINPUT45), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1018), .A2(KEYINPUT116), .A3(new_n1036), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1017), .A2(KEYINPUT116), .A3(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1016), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n499), .A2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1013), .A2(new_n1014), .B1(new_n1041), .B2(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1017), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1039), .A2(G1971), .B1(G2090), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G303), .A2(G8), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT55), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(G8), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n589), .A2(G1976), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT117), .B(G1976), .Z(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n714), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(G305), .B2(G1981), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n714), .A2(new_n1063), .A3(new_n1060), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1053), .B1(new_n1065), .B2(KEYINPUT49), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n1061), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1056), .B(new_n1059), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1044), .A2(KEYINPUT121), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1017), .B2(new_n1043), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1042), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n1039), .A2(G1971), .B1(new_n1073), .B2(G2090), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1049), .B1(new_n1074), .B2(G8), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1051), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1039), .A2(new_n804), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  INV_X1    g653(.A(G1961), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1077), .A2(new_n1078), .B1(new_n1079), .B2(new_n1045), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1018), .A2(new_n1036), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1078), .A2(G2078), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1015), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(G301), .B(KEYINPUT54), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(KEYINPUT125), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(KEYINPUT125), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1088), .A2(new_n1082), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1085), .B1(new_n1081), .B2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1084), .A2(new_n1085), .B1(new_n1080), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1015), .A2(new_n1018), .A3(new_n1036), .ZN(new_n1094));
  INV_X1    g669(.A(G1966), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G2084), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1042), .A2(new_n1097), .A3(new_n1044), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(G168), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1099), .B2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1093), .B1(new_n1101), .B2(G286), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1076), .B(new_n1092), .C1(new_n1100), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1015), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1073), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n840), .B(KEYINPUT57), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(KEYINPUT122), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1039), .A2(new_n1107), .B1(new_n1073), .B2(new_n1109), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1112), .B(KEYINPUT61), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1113), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(KEYINPUT124), .A3(KEYINPUT61), .A4(new_n1112), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1039), .A2(new_n1023), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n1129), .B2(new_n560), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1124), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n629), .B(new_n1131), .C1(new_n1125), .C2(new_n1128), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1130), .A2(new_n1132), .B1(KEYINPUT123), .B2(new_n1123), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1115), .A2(new_n1111), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1112), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1126), .A2(G2067), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1348), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n618), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n613), .B(new_n617), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(KEYINPUT60), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1122), .A2(new_n1133), .A3(new_n1137), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1120), .A2(new_n1142), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1112), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1105), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1074), .A2(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1048), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1126), .A2(G8), .A3(new_n1054), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT52), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1059), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1068), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1053), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1062), .ZN(new_n1157));
  NOR3_X1   g732(.A1(G305), .A2(KEYINPUT118), .A3(G1981), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1157), .A2(new_n1158), .B1(new_n1060), .B2(new_n714), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1159), .B2(new_n1067), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1154), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1052), .B(G286), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1151), .A2(new_n1161), .A3(new_n1050), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1046), .A2(G8), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1048), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1162), .A2(KEYINPUT63), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1161), .A4(new_n1050), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(G301), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT62), .B1(new_n1104), .B2(new_n1100), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1100), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1173), .B(new_n1174), .C1(new_n1103), .C2(new_n1102), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1076), .A2(new_n1171), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1053), .B(KEYINPUT119), .Z(new_n1177));
  NOR2_X1   g752(.A1(G288), .A2(G1976), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1064), .A2(new_n1062), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT120), .Z(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1051), .B2(new_n1161), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1170), .A2(new_n1176), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1035), .B1(new_n1149), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT48), .B1(new_n1034), .B2(new_n1019), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1034), .A2(KEYINPUT48), .A3(new_n1019), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1186), .B(new_n1187), .C1(new_n1019), .C2(new_n1029), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT46), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1026), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1019), .B1(new_n761), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT47), .Z(new_n1194));
  AND2_X1   g769(.A1(new_n1021), .A2(KEYINPUT126), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1028), .B1(new_n1021), .B2(KEYINPUT126), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1195), .A2(new_n1196), .B1(G2067), .B2(new_n791), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1188), .B(new_n1194), .C1(new_n1019), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g774(.A1(G229), .A2(new_n462), .A3(new_n664), .A4(G227), .ZN(new_n1201));
  AND2_X1   g775(.A1(new_n909), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n1202), .A2(new_n1004), .A3(new_n1002), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


