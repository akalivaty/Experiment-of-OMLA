//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n215), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  INV_X1    g0019(.A(new_n202), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT66), .B(G238), .Z(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G107), .A2(G264), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n209), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n212), .B(new_n223), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G232), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  OAI211_X1 g0050(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n252), .B1(new_n257), .B2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1698), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(G222), .B1(new_n266), .B2(G77), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n262), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n217), .A2(new_n253), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G169), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n207), .A2(G33), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT68), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n214), .A2(new_n216), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G50), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n281), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n206), .A2(G20), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n214), .A2(new_n216), .A3(new_n285), .A4(new_n282), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n287), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n275), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n294), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n272), .A2(G200), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n272), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n296), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(G226), .B(new_n308), .C1(new_n264), .C2(new_n265), .ZN(new_n309));
  OAI211_X1 g0109(.A(G232), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G97), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n217), .A2(new_n253), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n252), .B1(new_n257), .B2(G238), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT14), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(G169), .C1(new_n317), .C2(new_n318), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n317), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n225), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n279), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n283), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n332));
  INV_X1    g0132(.A(G13), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G1), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G20), .A3(new_n225), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n337));
  INV_X1    g0137(.A(new_n289), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n225), .B1(new_n206), .B2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n336), .A2(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n325), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G244), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n251), .B1(new_n256), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n268), .A2(G232), .A3(new_n308), .ZN(new_n345));
  INV_X1    g0145(.A(G107), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n268), .A2(G1698), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n345), .B1(new_n346), .B2(new_n268), .C1(new_n347), .C2(new_n224), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(new_n313), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G179), .ZN(new_n350));
  INV_X1    g0150(.A(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n349), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n353), .A2(new_n278), .B1(new_n207), .B2(new_n327), .ZN(new_n354));
  INV_X1    g0154(.A(new_n276), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n280), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n283), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n285), .A2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT70), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n338), .A2(G77), .A3(new_n288), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n318), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n301), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n317), .B2(new_n318), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n341), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n348), .A2(new_n313), .ZN(new_n371));
  INV_X1    g0171(.A(new_n344), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n361), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT71), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n349), .A2(G190), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n374), .A2(new_n376), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  AND4_X1   g0180(.A1(new_n342), .A2(new_n363), .A3(new_n370), .A4(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n266), .B2(new_n207), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n262), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G58), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n225), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n202), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n276), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n382), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n261), .A2(new_n207), .A3(new_n262), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n225), .B1(new_n396), .B2(new_n384), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n283), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n280), .A2(new_n286), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n292), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n290), .B1(new_n206), .B2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n280), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n251), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n407), .B2(new_n251), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(G223), .B(new_n308), .C1(new_n264), .C2(new_n265), .ZN(new_n413));
  OAI211_X1 g0213(.A(G226), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n313), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n351), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n407), .A2(new_n251), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT72), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n417), .A2(new_n420), .A3(G179), .A4(new_n409), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT73), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(new_n420), .A3(new_n409), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G169), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT73), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n421), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n406), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT18), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n406), .A2(new_n423), .A3(new_n430), .A4(new_n427), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT74), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n412), .A2(new_n433), .A3(new_n301), .A4(new_n417), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT74), .B1(new_n424), .B2(new_n367), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n424), .A2(G190), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n283), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT16), .B1(new_n397), .B2(new_n391), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n386), .A2(new_n382), .A3(new_n392), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n400), .B1(new_n293), .B2(new_n280), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT17), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n437), .A2(new_n443), .A3(KEYINPUT17), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n307), .A2(new_n381), .A3(new_n432), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT75), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT21), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT20), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  INV_X1    g0254(.A(G97), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n207), .C1(G33), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT83), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(new_n260), .B2(G97), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT83), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n283), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n453), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n456), .A2(new_n457), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(KEYINPUT20), .A3(new_n283), .A4(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n285), .A2(new_n462), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n260), .A2(G1), .ZN(new_n471));
  OAI21_X1  g0271(.A(G116), .B1(new_n289), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n465), .A2(new_n469), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G303), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G303), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n263), .A2(G257), .B1(new_n478), .B2(new_n266), .ZN(new_n479));
  OAI211_X1 g0279(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n271), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G41), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n206), .B(G45), .C1(new_n482), .C2(KEYINPUT5), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G41), .ZN(new_n485));
  OAI211_X1 g0285(.A(G270), .B(new_n254), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(G41), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(new_n206), .A3(G45), .A4(G274), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT79), .B1(new_n484), .B2(G41), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT79), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n482), .A3(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n486), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(G169), .B1(new_n481), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n452), .B1(new_n473), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n481), .A2(G190), .A3(new_n493), .ZN(new_n496));
  INV_X1    g0296(.A(new_n486), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n492), .A2(new_n488), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(new_n308), .C1(new_n264), .C2(new_n265), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT82), .B(G303), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n480), .B(new_n500), .C1(new_n268), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n313), .ZN(new_n503));
  AOI21_X1  g0303(.A(G200), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n473), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n351), .B1(new_n499), .B2(new_n503), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n493), .B1(new_n313), .B2(new_n502), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(KEYINPUT21), .B1(new_n507), .B2(G179), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n495), .B(new_n505), .C1(new_n473), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n289), .A2(new_n471), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n334), .A2(G20), .A3(new_n346), .ZN(new_n513));
  OR2_X1    g0313(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n207), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n268), .A2(new_n520), .A3(new_n207), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n346), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT23), .B1(new_n346), .B2(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n523), .A2(new_n524), .B1(G20), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(KEYINPUT24), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n283), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n519), .B2(new_n521), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(KEYINPUT24), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n511), .B(new_n517), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G264), .B(new_n254), .C1(new_n483), .C2(new_n485), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(new_n308), .C1(new_n264), .C2(new_n265), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n268), .A2(new_n537), .A3(G250), .A4(new_n308), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G294), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n536), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n534), .B1(new_n541), .B2(new_n313), .ZN(new_n542));
  INV_X1    g0342(.A(new_n498), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(G179), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n351), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n532), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n517), .A2(new_n511), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n530), .A2(KEYINPUT24), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n438), .B1(new_n530), .B2(KEYINPUT24), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(G200), .B1(new_n542), .B2(new_n543), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n539), .B(new_n540), .C1(new_n535), .C2(KEYINPUT85), .ZN(new_n552));
  INV_X1    g0352(.A(G250), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n261), .B2(new_n262), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n537), .B1(new_n554), .B2(new_n308), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n313), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  AND4_X1   g0356(.A1(new_n301), .A2(new_n556), .A3(new_n543), .A4(new_n533), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n550), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n546), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n285), .A2(G97), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT78), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(G97), .B2(new_n510), .ZN(new_n562));
  OAI21_X1  g0362(.A(G107), .B1(new_n383), .B2(new_n385), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n455), .A2(new_n346), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G97), .A2(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT6), .A2(G97), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(G107), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n346), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n276), .A2(G77), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n563), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n576), .A2(KEYINPUT77), .A3(new_n283), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT77), .B1(new_n576), .B2(new_n283), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n562), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n268), .A2(G250), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n308), .B1(new_n580), .B2(KEYINPUT4), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT4), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(G1698), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(G244), .C1(new_n265), .C2(new_n264), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n343), .B1(new_n261), .B2(new_n262), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n454), .C1(new_n585), .C2(KEYINPUT4), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n313), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G257), .B(new_n254), .C1(new_n483), .C2(new_n485), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n498), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G169), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n274), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n510), .A2(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n353), .A2(new_n286), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n207), .B1(new_n311), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G87), .A2(G97), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n346), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n207), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT80), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n597), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n283), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n598), .A2(new_n600), .B1(new_n597), .B2(new_n604), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n603), .B1(new_n608), .B2(new_n602), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n595), .B(new_n596), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(G238), .B(new_n308), .C1(new_n264), .C2(new_n265), .ZN(new_n611));
  OAI21_X1  g0411(.A(G244), .B1(new_n264), .B2(new_n265), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n525), .C1(new_n612), .C2(new_n308), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n313), .ZN(new_n614));
  INV_X1    g0414(.A(G45), .ZN(new_n615));
  OAI21_X1  g0415(.A(G250), .B1(new_n615), .B2(G1), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n254), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n367), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n613), .A2(new_n313), .B1(new_n254), .B2(new_n618), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n301), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n610), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n353), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n510), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n626), .B(new_n596), .C1(new_n607), .C2(new_n609), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT81), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT80), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n283), .A3(new_n606), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT81), .A3(new_n596), .A4(new_n626), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n622), .A2(G179), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n351), .B2(new_n622), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n624), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n587), .A2(new_n301), .A3(new_n590), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n543), .A2(new_n588), .ZN(new_n639));
  OAI21_X1  g0439(.A(G1698), .B1(new_n554), .B2(new_n582), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n612), .A2(new_n582), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n454), .A3(new_n584), .A4(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n313), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n638), .B1(new_n643), .B2(G200), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n644), .B(new_n562), .C1(new_n578), .C2(new_n577), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n594), .A2(new_n637), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n451), .A2(new_n509), .A3(new_n559), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n594), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n637), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n634), .A2(new_n636), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n646), .A2(new_n558), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n508), .A2(new_n473), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n465), .A2(new_n469), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n472), .A2(new_n470), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT21), .B1(new_n659), .B2(new_n506), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n655), .B1(new_n662), .B2(new_n546), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n450), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n305), .A2(new_n306), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n448), .A2(new_n370), .ZN(new_n667));
  INV_X1    g0467(.A(new_n341), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n319), .A2(KEYINPUT14), .B1(new_n323), .B2(G179), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n322), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n362), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n432), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n296), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n665), .A2(new_n673), .ZN(G369));
  INV_X1    g0474(.A(new_n546), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n334), .A2(new_n207), .ZN(new_n676));
  OAI21_X1  g0476(.A(G213), .B1(new_n676), .B2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT87), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT87), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(new_n680), .A3(KEYINPUT27), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n532), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n675), .B1(new_n558), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n546), .A2(new_n684), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n659), .A2(new_n684), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n509), .B2(KEYINPUT88), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n662), .A2(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT89), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(KEYINPUT90), .B(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n689), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n694), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n688), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n661), .A2(new_n684), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n687), .B1(new_n688), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT92), .Z(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  INV_X1    g0505(.A(new_n210), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(G41), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n210), .A2(KEYINPUT93), .A3(new_n482), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n206), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n599), .A2(new_n346), .A3(new_n462), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n711), .A2(new_n713), .B1(new_n222), .B2(new_n710), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  NAND2_X1  g0515(.A1(new_n664), .A2(new_n683), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n655), .B1(new_n661), .B2(new_n546), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n683), .B1(new_n654), .B2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(new_n717), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n559), .A2(new_n509), .A3(new_n684), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n622), .A2(new_n499), .A3(G179), .A4(new_n503), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n643), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n587), .A2(new_n533), .A3(new_n556), .A4(new_n590), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT94), .B(new_n728), .C1(new_n729), .C2(new_n725), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n542), .A2(new_n543), .ZN(new_n731));
  AOI21_X1  g0531(.A(G179), .B1(new_n499), .B2(new_n503), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n620), .A3(new_n591), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n481), .A2(new_n274), .A3(new_n493), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n643), .A3(new_n542), .A4(new_n622), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT94), .B1(new_n736), .B2(new_n728), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n684), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n724), .A2(new_n646), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n727), .A2(new_n733), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n736), .A2(new_n728), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT31), .B(new_n684), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n696), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n715), .B1(new_n745), .B2(G1), .ZN(G364));
  NOR2_X1   g0546(.A1(new_n698), .A2(new_n699), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n333), .A2(G20), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G45), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n711), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n747), .B(new_n750), .C1(new_n695), .C2(new_n697), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT95), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n207), .A2(new_n301), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n274), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n367), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G87), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n387), .A2(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n274), .A2(new_n367), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n207), .A2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n266), .B(new_n759), .C1(G68), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n207), .B1(new_n765), .B2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G97), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n761), .A2(new_n765), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n761), .A2(new_n754), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n756), .A2(new_n761), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n327), .A2(new_n773), .B1(new_n774), .B2(new_n346), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n753), .A2(new_n760), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G50), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n764), .A2(new_n768), .A3(new_n772), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(KEYINPUT33), .A2(G317), .ZN(new_n780));
  AND2_X1   g0580(.A1(KEYINPUT33), .A2(G317), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n763), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n774), .ZN(new_n784));
  INV_X1    g0584(.A(new_n769), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G329), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n755), .A2(new_n787), .B1(new_n773), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G294), .B2(new_n767), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n776), .B(KEYINPUT96), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT97), .B(G326), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n786), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n266), .B1(new_n757), .B2(new_n474), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  OAI21_X1  g0595(.A(new_n779), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n218), .B1(G20), .B2(new_n351), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n706), .A2(new_n266), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n462), .B2(new_n706), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n222), .A2(G45), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n246), .B2(G45), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n706), .A2(new_n268), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n797), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n750), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT99), .ZN(new_n812));
  INV_X1    g0612(.A(new_n808), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n695), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n752), .A2(new_n814), .ZN(G396));
  INV_X1    g0615(.A(new_n797), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n807), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G77), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT100), .B(G283), .Z(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n819), .A2(new_n762), .B1(new_n755), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n268), .B(new_n821), .C1(G303), .C2(new_n777), .ZN(new_n822));
  INV_X1    g0622(.A(new_n774), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G87), .A2(new_n823), .B1(new_n785), .B2(G311), .ZN(new_n824));
  INV_X1    g0624(.A(new_n757), .ZN(new_n825));
  INV_X1    g0625(.A(new_n773), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G107), .A2(new_n825), .B1(new_n826), .B2(G116), .ZN(new_n827));
  AND4_X1   g0627(.A1(new_n768), .A2(new_n822), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n777), .A2(G137), .B1(new_n826), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n755), .C1(new_n833), .C2(new_n762), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n835));
  XNOR2_X1  g0635(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n268), .B1(new_n757), .B2(new_n284), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n774), .A2(new_n225), .B1(new_n769), .B2(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n837), .B(new_n839), .C1(G58), .C2(new_n767), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n830), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n750), .B(new_n818), .C1(new_n843), .C2(new_n797), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n377), .A2(new_n683), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n380), .A2(new_n846), .B1(new_n361), .B2(new_n352), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n352), .A2(new_n361), .A3(new_n683), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT103), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n349), .A2(G190), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n349), .A2(new_n367), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n378), .A2(new_n376), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n845), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n851), .B(new_n848), .C1(new_n856), .C2(new_n362), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n844), .B1(new_n859), .B2(new_n807), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n716), .B(new_n859), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n744), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n750), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n861), .A2(new_n744), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(G384));
  XOR2_X1   g0665(.A(new_n573), .B(KEYINPUT104), .Z(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT35), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(KEYINPUT35), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(G116), .A3(new_n219), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OR3_X1    g0670(.A1(new_n221), .A2(new_n327), .A3(new_n388), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n201), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n206), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT111), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n451), .B2(new_n722), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n723), .A2(KEYINPUT111), .A3(new_n450), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n876), .A2(new_n877), .A3(new_n673), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n664), .A2(new_n683), .A3(new_n859), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n879), .A2(new_n848), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n668), .A2(new_n683), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT105), .B1(new_n342), .B2(new_n370), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT105), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n883), .B(new_n369), .C1(new_n325), .C2(new_n341), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n670), .B2(new_n369), .ZN(new_n886));
  INV_X1    g0686(.A(new_n881), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n342), .A2(KEYINPUT105), .A3(new_n370), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n429), .A2(new_n446), .A3(new_n431), .A4(new_n447), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n406), .A2(new_n682), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n427), .B1(new_n441), .B2(new_n442), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n426), .B1(new_n425), .B2(new_n421), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT106), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n406), .A2(new_n423), .A3(new_n900), .A4(new_n427), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n682), .B(KEYINPUT107), .Z(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT37), .B1(new_n406), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n899), .A2(new_n444), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n428), .A2(new_n444), .A3(new_n894), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n896), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT108), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(KEYINPUT108), .A3(new_n911), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n892), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n896), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n896), .B2(new_n907), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT39), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n406), .A2(new_n902), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n428), .A2(new_n444), .A3(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n893), .A2(new_n920), .B1(new_n904), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT109), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n911), .A2(KEYINPUT110), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n893), .A2(new_n920), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n904), .A2(new_n922), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT109), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n909), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT110), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n896), .A2(new_n907), .A3(new_n931), .A4(KEYINPUT38), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n924), .A2(new_n925), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n918), .B1(new_n933), .B2(KEYINPUT39), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n342), .A2(new_n684), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n432), .A2(new_n902), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n915), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n878), .B(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n738), .A2(new_n739), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n451), .B1(new_n740), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n933), .A2(KEYINPUT40), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n858), .B1(new_n740), .B2(new_n940), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT113), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n943), .A2(new_n944), .A3(new_n890), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n943), .B2(new_n890), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n890), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n916), .B2(new_n917), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n950), .B2(new_n913), .ZN(new_n951));
  XNOR2_X1  g0751(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n942), .A2(new_n947), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n941), .B(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n696), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n939), .A2(new_n957), .B1(new_n206), .B2(new_n748), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n939), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n874), .B1(new_n958), .B2(new_n959), .ZN(G367));
  OAI21_X1  g0760(.A(new_n809), .B1(new_n210), .B2(new_n353), .ZN(new_n961));
  INV_X1    g0761(.A(new_n242), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n803), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n750), .A2(new_n963), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n819), .A2(new_n773), .B1(new_n755), .B2(new_n501), .ZN(new_n965));
  INV_X1    g0765(.A(G317), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n762), .A2(new_n820), .B1(new_n769), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n791), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n965), .B(new_n967), .C1(new_n968), .C2(G311), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n825), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n268), .B1(new_n823), .B2(G97), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT46), .B1(new_n825), .B2(G116), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G107), .B2(new_n767), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n823), .A2(G77), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n770), .B2(new_n762), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n766), .A2(new_n225), .ZN(new_n977));
  INV_X1    g0777(.A(G137), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n268), .B1(new_n769), .B2(new_n978), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n201), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n826), .A2(new_n981), .B1(new_n825), .B2(G58), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n833), .B2(new_n755), .C1(new_n791), .C2(new_n832), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n974), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n797), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(new_n637), .ZN(new_n989));
  INV_X1    g0789(.A(new_n610), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(new_n990), .B2(new_n683), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n652), .A2(new_n610), .A3(new_n684), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n964), .B1(new_n987), .B2(new_n988), .C1(new_n994), .C2(new_n813), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n749), .A2(G1), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n747), .B1(new_n687), .B2(new_n686), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n700), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n661), .B2(new_n684), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n700), .A3(new_n701), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n579), .A2(new_n684), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n594), .A2(new_n1002), .A3(new_n645), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n594), .B2(new_n683), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n703), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT44), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n703), .A2(new_n1004), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n700), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n745), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n709), .B(KEYINPUT41), .Z(new_n1014));
  AOI21_X1  g0814(.A(new_n996), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1004), .B(KEYINPUT114), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n675), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n684), .B1(new_n1019), .B2(new_n594), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n688), .A2(new_n701), .A3(new_n1004), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT42), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1018), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1017), .B(new_n1025), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n995), .B1(new_n1015), .B2(new_n1027), .ZN(G387));
  NAND3_X1  g0828(.A1(new_n999), .A2(new_n745), .A3(new_n1000), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n710), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n745), .B1(new_n999), .B2(new_n1000), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n999), .A2(new_n1000), .A3(new_n996), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n238), .A2(G45), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n404), .A2(new_n284), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n713), .B(new_n615), .C1(new_n225), .C2(new_n327), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1035), .B(new_n803), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n799), .A2(new_n712), .B1(new_n346), .B2(new_n706), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n750), .B1(new_n1041), .B2(new_n809), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n755), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G50), .A2(new_n1043), .B1(new_n785), .B2(G150), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n268), .C1(new_n455), .C2(new_n774), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n762), .A2(new_n280), .B1(new_n773), .B2(new_n225), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n776), .A2(new_n770), .B1(new_n757), .B2(new_n327), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n766), .A2(new_n353), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n266), .B1(new_n769), .B2(new_n792), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G317), .A2(new_n1043), .B1(new_n826), .B2(new_n478), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n788), .B2(new_n762), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G322), .B2(new_n968), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1053), .A2(KEYINPUT48), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n819), .A2(new_n766), .B1(new_n757), .B2(new_n820), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(KEYINPUT48), .B2(new_n1053), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1050), .B(new_n1059), .C1(G116), .C2(new_n823), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1049), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1042), .B1(new_n688), .B2(new_n813), .C1(new_n1062), .C2(new_n816), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT117), .Z(new_n1064));
  NAND2_X1  g0864(.A1(new_n1034), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1033), .A2(new_n1066), .ZN(G393));
  INV_X1    g0867(.A(new_n1029), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1012), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n709), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1016), .A2(new_n813), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n776), .A2(new_n833), .B1(new_n755), .B2(new_n770), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n268), .B1(new_n766), .B2(new_n327), .C1(new_n758), .C2(new_n774), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n757), .A2(new_n225), .B1(new_n769), .B2(new_n832), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n201), .A2(new_n762), .B1(new_n773), .B2(new_n280), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n776), .A2(new_n966), .B1(new_n755), .B2(new_n788), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n266), .B1(new_n766), .B2(new_n462), .C1(new_n346), .C2(new_n774), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n762), .A2(new_n501), .B1(new_n769), .B2(new_n787), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n819), .A2(new_n757), .B1(new_n773), .B2(new_n820), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1074), .A2(new_n1078), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(new_n816), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n809), .B1(new_n455), .B2(new_n210), .C1(new_n804), .C2(new_n249), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n750), .B1(new_n1087), .B2(KEYINPUT118), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(KEYINPUT118), .B2(new_n1087), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1072), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1069), .B2(new_n996), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1071), .A2(new_n1091), .ZN(G390));
  NAND2_X1  g0892(.A1(new_n941), .A2(G330), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1093), .A2(new_n876), .A3(new_n673), .A4(new_n877), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n943), .A2(G330), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n891), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n744), .A2(new_n859), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n891), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n880), .A2(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n720), .A2(new_n858), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(new_n848), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1095), .A2(new_n891), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n744), .A2(new_n890), .A3(new_n859), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1099), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1094), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n933), .B1(new_n342), .B2(new_n684), .C1(new_n1101), .C2(new_n891), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n892), .A2(new_n935), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n934), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1096), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1108), .B(new_n1103), .C1(new_n1109), .C2(new_n934), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n709), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1106), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n750), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n823), .A2(new_n981), .B1(new_n763), .B2(G137), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n769), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT53), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n757), .B2(new_n833), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n825), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n268), .B1(new_n755), .B2(new_n838), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n776), .A2(new_n1126), .B1(new_n773), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1125), .B(new_n1128), .C1(G159), .C2(new_n767), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n266), .B1(new_n757), .B2(new_n758), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n225), .A2(new_n774), .B1(new_n773), .B2(new_n455), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(G77), .C2(new_n767), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n776), .A2(new_n783), .B1(new_n762), .B2(new_n346), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n755), .A2(new_n462), .B1(new_n769), .B2(new_n820), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1124), .A2(new_n1129), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1117), .B1(new_n404), .B2(new_n817), .C1(new_n1136), .C2(new_n816), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT119), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n934), .B2(new_n807), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n996), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1113), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1116), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G378));
  OAI21_X1  g0943(.A(new_n1117), .B1(new_n981), .B2(new_n817), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n755), .A2(new_n346), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT120), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n777), .A2(G116), .B1(new_n826), .B2(new_n625), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n783), .C2(new_n769), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n482), .B(new_n266), .C1(new_n757), .C2(new_n327), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n762), .A2(new_n455), .B1(new_n774), .B2(new_n387), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1148), .A2(new_n977), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n266), .A2(new_n482), .ZN(new_n1152));
  AOI21_X1  g0952(.A(G50), .B1(new_n260), .B2(new_n482), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1151), .A2(KEYINPUT58), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n776), .A2(new_n1119), .B1(new_n762), .B2(new_n838), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n826), .A2(G137), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n1126), .B2(new_n755), .C1(new_n757), .C2(new_n1127), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G150), .C2(new_n767), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n260), .B(new_n482), .C1(new_n774), .C2(new_n770), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G124), .B2(new_n785), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT59), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1154), .B1(KEYINPUT58), .B2(new_n1151), .C1(new_n1160), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1144), .B1(new_n1165), .B2(new_n797), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n294), .A2(new_n682), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n307), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n307), .A2(new_n1167), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  OR3_X1    g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1166), .B1(new_n1173), .B2(new_n807), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n955), .A2(new_n1173), .A3(G330), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  INV_X1    g0977(.A(G330), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n954), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n948), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n914), .B2(new_n912), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n952), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n933), .B(KEYINPUT40), .C1(new_n945), .C2(new_n946), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1182), .A2(KEYINPUT121), .A3(G330), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1173), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT122), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT122), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1188), .B(new_n1173), .C1(new_n1179), .C2(new_n1184), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1176), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n938), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n938), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1176), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1175), .B1(new_n1194), .B2(new_n996), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1115), .A2(new_n878), .A3(new_n1093), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1196), .A2(new_n1194), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n710), .B1(new_n1197), .B2(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1188), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1185), .A2(KEYINPUT122), .A3(new_n1186), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1202), .A2(KEYINPUT123), .A3(new_n1192), .A4(new_n1176), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT123), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1193), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1205), .A3(new_n1191), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1196), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1195), .B1(new_n1198), .B2(new_n1207), .ZN(G375));
  NAND2_X1  g1008(.A1(new_n1094), .A2(new_n1105), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1107), .A2(new_n1014), .A3(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1105), .A2(new_n1140), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1117), .B1(G68), .B2(new_n817), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G150), .A2(new_n826), .B1(new_n785), .B2(G128), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n770), .B2(new_n757), .C1(new_n762), .C2(new_n1127), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G132), .A2(new_n777), .B1(new_n1043), .B2(G137), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n266), .B1(new_n823), .B2(G58), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n284), .C2(new_n766), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n825), .B1(new_n785), .B2(G303), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n346), .B2(new_n773), .C1(new_n820), .C2(new_n776), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G116), .A2(new_n763), .B1(new_n1043), .B2(G283), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1048), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1220), .A2(new_n266), .A3(new_n975), .A4(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1214), .A2(new_n1217), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1212), .B1(new_n797), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n890), .B2(new_n807), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1210), .A2(new_n1211), .A3(new_n1225), .ZN(G381));
  OR2_X1    g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G387), .ZN(new_n1229));
  INV_X1    g1029(.A(G396), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1033), .A2(new_n1230), .A3(new_n1066), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(G390), .A2(new_n1231), .A3(G384), .A4(G381), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1229), .A3(new_n1232), .ZN(G407));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1227), .ZN(G409));
  OAI21_X1  g1034(.A(G396), .B1(new_n1032), .B2(new_n1065), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1229), .B2(KEYINPUT127), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G387), .A2(new_n1231), .A3(new_n1235), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1237), .A2(G390), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G390), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G213), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(G343), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1175), .B1(new_n1206), .B2(new_n996), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(KEYINPUT124), .B(new_n1175), .C1(new_n1206), .C2(new_n996), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1196), .A2(new_n1014), .A3(new_n1194), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT125), .B1(new_n1251), .B2(new_n1142), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1253));
  OAI211_X1 g1053(.A(KEYINPUT125), .B(new_n1142), .C1(new_n1253), .C2(new_n1248), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1195), .C1(new_n1198), .C2(new_n1207), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1244), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1211), .A2(new_n1225), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1209), .B(KEYINPUT60), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1106), .A2(new_n709), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(G384), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1243), .A2(G2897), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1262), .B(new_n1263), .ZN(new_n1264));
  AOI211_X1 g1064(.A(KEYINPUT61), .B(new_n1241), .C1(new_n1257), .C2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1262), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1244), .B(new_n1266), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT63), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1265), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1142), .B1(new_n1253), .B2(new_n1248), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1243), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1264), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1267), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(KEYINPUT62), .A3(new_n1266), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1281), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1241), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1273), .B1(new_n1285), .B2(new_n1286), .ZN(G405));
  XNOR2_X1  g1087(.A(new_n1241), .B(new_n1262), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G375), .B(G378), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1288), .B(new_n1289), .ZN(G402));
endmodule


