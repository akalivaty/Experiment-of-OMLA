//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  XOR2_X1   g003(.A(G125), .B(G140), .Z(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(new_n187), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(KEYINPUT23), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n196), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G110), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n193), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n191), .A2(new_n192), .ZN(new_n204));
  XNOR2_X1  g018(.A(G125), .B(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n192), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n201), .A2(G110), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n204), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G137), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(KEYINPUT70), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n214));
  XOR2_X1   g028(.A(new_n212), .B(new_n214), .Z(new_n215));
  XNOR2_X1  g029(.A(new_n210), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G902), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G217), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G234), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n219), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n222), .A2(G902), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT31), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n192), .A2(G143), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n197), .A2(new_n192), .A3(G143), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n231), .B(G146), .C1(new_n197), .C2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(G134), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n247), .A3(G131), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT0), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(new_n197), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT0), .B(G128), .Z(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT65), .A2(G131), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n240), .A2(new_n243), .A3(new_n256), .A4(new_n241), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT66), .B1(new_n258), .B2(new_n259), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n263), .A3(KEYINPUT30), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n259), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n265), .A2(new_n255), .B1(new_n249), .B2(new_n236), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(G116), .B(G119), .Z(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT2), .B(G113), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n264), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n262), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n260), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n274), .A2(new_n255), .B1(new_n237), .B2(new_n249), .ZN(new_n275));
  INV_X1    g089(.A(new_n271), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G101), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n213), .A3(G210), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n272), .A2(new_n285), .A3(new_n277), .A4(new_n282), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n228), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n272), .A2(new_n277), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n228), .A3(new_n282), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n266), .A2(new_n276), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n277), .A2(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n277), .A2(KEYINPUT28), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n292), .B1(new_n296), .B2(new_n282), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI211_X1 g112(.A(KEYINPUT69), .B(new_n228), .C1(new_n284), .C2(new_n286), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n290), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n289), .A2(new_n299), .A3(new_n297), .ZN(new_n305));
  INV_X1    g119(.A(new_n303), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT32), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n291), .A2(new_n282), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT29), .B(new_n309), .C1(new_n296), .C2(new_n282), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n275), .A2(new_n276), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n294), .B2(new_n295), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT29), .A3(new_n282), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n217), .ZN(new_n314));
  OAI21_X1  g128(.A(G472), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n227), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G221), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT9), .B(G234), .Z(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(new_n217), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT3), .A2(G107), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT3), .A2(G107), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(G104), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  INV_X1    g137(.A(G107), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT71), .A2(G104), .ZN(new_n326));
  NOR2_X1   g140(.A1(KEYINPUT71), .A2(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(G104), .A2(G107), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(G101), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n236), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n236), .A3(new_n333), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT74), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n274), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n342), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n338), .A2(KEYINPUT12), .A3(new_n265), .A4(new_n340), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OR2_X1    g162(.A1(KEYINPUT71), .A2(G104), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT71), .A2(G104), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n321), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT3), .A2(G107), .ZN(new_n352));
  INV_X1    g166(.A(G104), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n325), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n330), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n355), .A2(KEYINPUT72), .A3(KEYINPUT4), .A4(new_n330), .ZN(new_n359));
  INV_X1    g173(.A(new_n355), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n358), .A2(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n255), .ZN(new_n363));
  INV_X1    g177(.A(new_n274), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n337), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n237), .A2(KEYINPUT10), .A3(new_n330), .A4(new_n333), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(new_n364), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G140), .ZN(new_n369));
  INV_X1    g183(.A(G227), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G953), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n369), .B(new_n371), .Z(new_n372));
  NAND3_X1  g186(.A1(new_n348), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n274), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n368), .ZN(new_n377));
  INV_X1    g191(.A(new_n372), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n348), .A2(new_n380), .A3(new_n368), .A4(new_n372), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n217), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n382), .A2(KEYINPUT77), .A3(new_n383), .A4(new_n217), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n348), .A2(new_n368), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n378), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n368), .A3(new_n372), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n217), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G469), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n319), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(G214), .B1(G237), .B2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n358), .A2(new_n359), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n360), .A2(new_n361), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n271), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT78), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n195), .A3(G116), .ZN(new_n404));
  OAI211_X1 g218(.A(G113), .B(new_n404), .C1(new_n269), .C2(new_n403), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n269), .B2(new_n270), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n406), .A2(new_n334), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n362), .A2(new_n408), .A3(new_n271), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n398), .B1(new_n413), .B2(KEYINPUT6), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n415), .A4(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n410), .A2(new_n412), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n419));
  INV_X1    g233(.A(new_n255), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G125), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(G125), .B2(new_n236), .ZN(new_n422));
  MUX2_X1   g236(.A(new_n421), .B(new_n422), .S(KEYINPUT81), .Z(new_n423));
  NAND2_X1  g237(.A1(new_n213), .A2(G224), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT82), .Z(new_n425));
  XOR2_X1   g239(.A(new_n423), .B(new_n425), .Z(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(KEYINPUT7), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n423), .A2(new_n428), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n406), .A2(new_n334), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n407), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n412), .B(KEYINPUT8), .Z(new_n434));
  NAND3_X1  g248(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n334), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n418), .A2(new_n429), .A3(new_n430), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n427), .A2(new_n217), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n427), .A2(new_n217), .A3(new_n439), .A4(new_n437), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n397), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G475), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n280), .A2(new_n213), .A3(G214), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(G143), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n245), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT18), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n446), .B1(new_n449), .B2(new_n245), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n190), .A2(G146), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n206), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(KEYINPUT17), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n446), .B(new_n245), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(KEYINPUT17), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n456), .B2(new_n193), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n353), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT19), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n455), .B(new_n204), .C1(G146), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n459), .B1(new_n464), .B2(new_n453), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n444), .B(new_n217), .C1(new_n461), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n460), .B2(new_n457), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n444), .A4(new_n217), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n471), .A3(KEYINPUT20), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n457), .B(new_n459), .ZN(new_n473));
  OAI21_X1  g287(.A(G475), .B1(new_n473), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n466), .A2(KEYINPUT85), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G952), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT21), .B(G898), .Z(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n486));
  AND2_X1   g300(.A1(KEYINPUT86), .A2(G122), .ZN(new_n487));
  NOR2_X1   g301(.A1(KEYINPUT86), .A2(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(G116), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT87), .Z(new_n490));
  INV_X1    g304(.A(G116), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G122), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(KEYINPUT14), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(G107), .ZN(new_n495));
  XNOR2_X1  g309(.A(G128), .B(G143), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n239), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n490), .B(new_n492), .C1(KEYINPUT14), .C2(new_n324), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(KEYINPUT13), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n197), .A2(KEYINPUT13), .A3(G143), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n239), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n500), .A2(new_n502), .B1(new_n239), .B2(new_n496), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n490), .A2(new_n324), .A3(new_n492), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n324), .B1(new_n490), .B2(new_n492), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n318), .A2(G217), .A3(new_n213), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n510));
  INV_X1    g324(.A(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n499), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n499), .A2(KEYINPUT88), .A3(new_n506), .A4(new_n511), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n217), .A4(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G478), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n516), .A2(new_n518), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n486), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n516), .A2(new_n518), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT90), .A3(new_n519), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n477), .B(new_n485), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n316), .A2(new_n395), .A3(new_n443), .A4(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT91), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(G3));
  INV_X1    g342(.A(G472), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n301), .B2(new_n217), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(KEYINPUT92), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n532));
  OAI21_X1  g346(.A(G472), .B1(new_n305), .B2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n301), .A2(new_n303), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n227), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n397), .B(new_n485), .C1(new_n441), .C2(new_n442), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n536), .A2(new_n395), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n513), .A2(new_n217), .A3(new_n515), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n513), .A2(new_n542), .A3(new_n515), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n507), .B2(new_n508), .ZN(new_n545));
  AOI211_X1 g359(.A(KEYINPUT93), .B(new_n511), .C1(new_n499), .C2(new_n506), .ZN(new_n546));
  OAI211_X1 g360(.A(KEYINPUT33), .B(new_n512), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n547), .A3(new_n217), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n541), .B1(new_n548), .B2(new_n517), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n477), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT94), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n539), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT34), .B(G104), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(G6));
  AND2_X1   g368(.A1(new_n522), .A2(new_n524), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n539), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT35), .B(G107), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(G9));
  NAND3_X1  g374(.A1(new_n395), .A2(new_n443), .A3(new_n525), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n215), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n566), .B(new_n210), .Z(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n225), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n224), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT97), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n536), .A3(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(G110), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n571), .B(new_n573), .ZN(G12));
  NAND2_X1  g388(.A1(new_n308), .A2(new_n315), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n395), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n441), .A2(new_n442), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n396), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n481), .B(KEYINPUT99), .Z(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(G900), .B2(new_n483), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT100), .Z(new_n585));
  NOR2_X1   g399(.A1(new_n557), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n577), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT101), .B(G128), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G30));
  NAND2_X1  g403(.A1(new_n284), .A2(new_n286), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n311), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n282), .B1(new_n592), .B2(new_n277), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n217), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G472), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n569), .B1(new_n308), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n585), .B(KEYINPUT102), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(KEYINPUT39), .Z(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n395), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(KEYINPUT40), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n601), .A2(KEYINPUT40), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n579), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n522), .A2(new_n524), .A3(new_n477), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n441), .A2(KEYINPUT38), .A3(new_n442), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n602), .A2(new_n603), .A3(new_n396), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G143), .ZN(G45));
  NOR2_X1   g424(.A1(new_n550), .A2(new_n585), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n577), .A2(new_n581), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G146), .ZN(G48));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n614));
  INV_X1    g428(.A(new_n319), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n383), .B1(new_n382), .B2(new_n217), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AND4_X1   g431(.A1(new_n614), .A2(new_n388), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n386), .B2(new_n387), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n614), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n316), .A3(new_n538), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n551), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT41), .B(G113), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G15));
  INV_X1    g439(.A(new_n557), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n621), .A2(new_n316), .A3(new_n538), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G116), .ZN(G18));
  NAND3_X1  g442(.A1(new_n388), .A2(new_n615), .A3(new_n617), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT103), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n619), .A2(new_n614), .A3(new_n615), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n443), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT104), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n630), .A2(new_n634), .A3(new_n443), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n525), .A3(new_n577), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G119), .ZN(G21));
  INV_X1    g452(.A(new_n606), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n303), .B(KEYINPUT105), .Z(new_n640));
  OAI21_X1  g454(.A(new_n292), .B1(new_n312), .B2(new_n282), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n287), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n533), .A3(new_n537), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n621), .A2(new_n538), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G122), .ZN(G24));
  NAND3_X1  g462(.A1(new_n644), .A2(new_n533), .A3(new_n569), .ZN(new_n649));
  INV_X1    g463(.A(new_n611), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n634), .B1(new_n621), .B2(new_n443), .ZN(new_n652));
  INV_X1    g466(.A(new_n635), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G125), .ZN(G27));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n390), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n389), .A2(KEYINPUT107), .A3(new_n378), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n391), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n383), .B1(new_n659), .B2(new_n217), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n388), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n615), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n386), .B2(new_n387), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT108), .B1(new_n665), .B2(new_n319), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n441), .A2(new_n396), .A3(new_n442), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(KEYINPUT42), .A3(new_n316), .A4(new_n611), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n316), .A2(new_n664), .A3(new_n666), .A4(new_n668), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n671), .B1(new_n672), .B2(new_n650), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G131), .ZN(G33));
  AND2_X1   g489(.A1(new_n586), .A2(KEYINPUT109), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n586), .A2(KEYINPUT109), .ZN(new_n677));
  OR3_X1    g491(.A1(new_n676), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G134), .ZN(G36));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n392), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g495(.A(G469), .B(new_n681), .C1(new_n659), .C2(new_n680), .ZN(new_n682));
  NAND2_X1  g496(.A1(G469), .A2(G902), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n682), .A2(KEYINPUT46), .A3(new_n683), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n388), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n615), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n599), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n556), .A2(new_n549), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n556), .A2(new_n549), .A3(KEYINPUT43), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n569), .B(new_n695), .C1(new_n535), .C2(new_n531), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n667), .B(new_n700), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n690), .A2(new_n698), .A3(new_n699), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n242), .ZN(G39));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n689), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n688), .A2(KEYINPUT47), .A3(new_n615), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n650), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n575), .A2(new_n537), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n668), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G140), .ZN(G42));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n715));
  INV_X1    g529(.A(new_n525), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n716), .B(new_n576), .C1(new_n633), .C2(new_n635), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n443), .A2(new_n484), .A3(new_n537), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n523), .A2(new_n519), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n556), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(new_n395), .A3(new_n536), .A4(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n627), .A2(new_n571), .A3(new_n647), .A4(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n717), .A2(new_n724), .A3(new_n623), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n305), .A2(new_n306), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT92), .B1(new_n530), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n533), .A2(new_n532), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n395), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n718), .A3(new_n550), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n575), .A2(new_n537), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n561), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n726), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(KEYINPUT112), .B(new_n526), .C1(new_n539), .C2(new_n550), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n674), .A2(new_n678), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n651), .A2(new_n664), .A3(new_n666), .A4(new_n668), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT113), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n578), .A2(new_n720), .A3(new_n585), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n577), .A3(new_n556), .A4(new_n668), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n725), .A2(new_n736), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n587), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n665), .A2(new_n319), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n596), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n585), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n443), .A2(new_n748), .A3(new_n606), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n745), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n749), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(KEYINPUT114), .A3(new_n596), .A4(new_n746), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n654), .A2(new_n744), .A3(new_n612), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT52), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n587), .B1(new_n636), .B2(new_n651), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n612), .A4(new_n753), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n715), .B1(new_n743), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n724), .ZN(new_n761));
  INV_X1    g575(.A(new_n623), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n736), .A3(new_n762), .A4(new_n637), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n674), .A2(new_n739), .A3(new_n678), .A4(new_n741), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT53), .A3(new_n755), .A4(new_n758), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n760), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(new_n760), .B2(new_n766), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n583), .B1(new_n693), .B2(new_n694), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n630), .A2(new_n772), .A3(new_n668), .A4(new_n631), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n732), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT48), .Z(new_n775));
  INV_X1    g589(.A(new_n645), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n772), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n636), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n773), .A2(new_n649), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n308), .A2(new_n595), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n630), .A3(new_n631), .A4(new_n668), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n227), .A2(new_n481), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n549), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n779), .B1(new_n784), .B2(new_n556), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n619), .A2(KEYINPUT116), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n619), .A2(KEYINPUT116), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n319), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n705), .A2(new_n706), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n777), .A2(new_n701), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n777), .A2(new_n701), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n396), .B1(new_n605), .B2(new_n607), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n777), .A2(new_n621), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n801), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n777), .A2(new_n621), .A3(new_n803), .A4(new_n798), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n785), .A2(new_n794), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n795), .A2(new_n796), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n778), .B(new_n479), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n782), .A2(new_n551), .A3(new_n783), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n771), .A2(KEYINPUT119), .A3(new_n775), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n760), .A2(new_n766), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT54), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n775), .A3(new_n812), .A4(new_n768), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n478), .A2(new_n213), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n619), .B(KEYINPUT49), .Z(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n227), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n319), .B1(new_n605), .B2(new_n607), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n780), .A2(new_n691), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n396), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n820), .A2(new_n825), .ZN(G75));
  AOI21_X1  g640(.A(new_n217), .B1(new_n760), .B2(new_n766), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT56), .B1(new_n827), .B2(G210), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n417), .A2(new_n419), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(new_n426), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT55), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n213), .A2(G952), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(G210), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n831), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n832), .A2(new_n834), .A3(new_n837), .ZN(G51));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n815), .A2(new_n839), .A3(new_n768), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n770), .A2(KEYINPUT120), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n683), .B(KEYINPUT57), .Z(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n382), .ZN(new_n844));
  INV_X1    g658(.A(new_n682), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n827), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n833), .B1(new_n844), .B2(new_n846), .ZN(G54));
  NAND3_X1  g661(.A1(new_n827), .A2(KEYINPUT58), .A3(G475), .ZN(new_n848));
  INV_X1    g662(.A(new_n469), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n851), .A3(new_n833), .ZN(G60));
  NAND2_X1  g666(.A1(new_n543), .A2(new_n547), .ZN(new_n853));
  NAND2_X1  g667(.A1(G478), .A2(G902), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT59), .Z(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n771), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n853), .A2(new_n855), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n840), .A2(new_n841), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n856), .A2(new_n858), .A3(new_n834), .ZN(G63));
  XNOR2_X1  g673(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n221), .A2(new_n217), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n814), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n567), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n834), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n863), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n216), .B(KEYINPUT122), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n866), .B(KEYINPUT61), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n865), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(G66));
  NAND2_X1  g687(.A1(new_n482), .A2(G224), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(G953), .ZN(new_n875));
  INV_X1    g689(.A(new_n763), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(G953), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT123), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n829), .B1(G898), .B2(new_n213), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(G69));
  AOI21_X1  g694(.A(new_n702), .B1(new_n711), .B2(new_n712), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n690), .A2(new_n443), .A3(new_n316), .A4(new_n606), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n612), .A3(new_n756), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n737), .A2(new_n213), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n883), .A2(new_n884), .B1(new_n370), .B2(new_n213), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n264), .A2(new_n268), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT124), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n463), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(G900), .B1(new_n888), .B2(G227), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(G953), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n654), .A2(new_n609), .A3(new_n744), .A4(new_n612), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n601), .A2(new_n667), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n721), .A2(new_n550), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n316), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n881), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT125), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n894), .A2(new_n881), .A3(new_n900), .A4(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n213), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n889), .B(new_n891), .C1(new_n903), .C2(new_n888), .ZN(G72));
  NAND2_X1  g718(.A1(G472), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT63), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n876), .A2(new_n737), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n883), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n282), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n909), .A3(new_n291), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n906), .B1(new_n591), .B2(new_n309), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n814), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n910), .A2(new_n834), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n899), .A2(new_n876), .A3(new_n901), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(KEYINPUT126), .A3(new_n906), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(new_n282), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT126), .B1(new_n917), .B2(new_n906), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n291), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n919), .B2(new_n921), .ZN(G57));
endmodule


