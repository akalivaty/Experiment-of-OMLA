//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AOI21_X1  g057(.A(new_n479), .B1(new_n469), .B2(new_n470), .ZN(new_n483));
  MUX2_X1   g058(.A(G100), .B(G112), .S(G2105), .Z(new_n484));
  AOI22_X1  g059(.A1(G124), .A2(new_n483), .B1(new_n484), .B2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n479), .B1(new_n463), .B2(new_n464), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT69), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n492), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT70), .B1(new_n492), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(new_n479), .C1(new_n464), .C2(new_n463), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n477), .A2(new_n502), .A3(new_n479), .A4(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(G651), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n510), .A2(G543), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT73), .B1(new_n515), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT5), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(new_n519), .B1(new_n515), .B2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n508), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(G166));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(new_n511), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n520), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n532));
  AND3_X1   g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n512), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n510), .A2(G543), .A3(new_n511), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n535), .B1(G51), .B2(new_n540), .ZN(G168));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n537), .B2(new_n539), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT76), .B(G90), .Z(new_n545));
  AOI22_X1  g120(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n521), .A2(new_n545), .B1(new_n546), .B2(new_n508), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n508), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n515), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n517), .B1(KEYINPUT5), .B2(new_n518), .ZN(new_n556));
  NOR3_X1   g131(.A1(new_n515), .A2(KEYINPUT73), .A3(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n560), .A2(KEYINPUT77), .A3(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n539), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n564));
  OAI21_X1  g139(.A(G43), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n528), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G81), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n514), .A2(new_n576), .A3(new_n520), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT78), .B1(new_n528), .B2(new_n558), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(new_n578), .A3(G91), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n508), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n510), .A2(G53), .A3(G543), .A4(new_n511), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT9), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  NAND3_X1  g161(.A1(new_n577), .A2(new_n578), .A3(G87), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n558), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(G651), .A2(new_n589), .B1(new_n512), .B2(G49), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT79), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n587), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G288));
  NAND3_X1  g171(.A1(new_n577), .A2(new_n578), .A3(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n558), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G48), .B2(new_n512), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n508), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(G85), .B2(new_n566), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n540), .A2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT80), .Z(new_n609));
  NAND3_X1  g184(.A1(new_n577), .A2(new_n578), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT10), .A4(G92), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n558), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n612), .A2(new_n613), .B1(G651), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n540), .A2(KEYINPUT81), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n537), .B2(new_n539), .ZN(new_n620));
  OAI21_X1  g195(.A(G54), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(G868), .B2(new_n623), .ZN(G284));
  OAI21_X1  g199(.A(new_n609), .B1(G868), .B2(new_n623), .ZN(G321));
  NOR2_X1   g200(.A1(G299), .A2(G868), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g202(.A(new_n626), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND3_X1  g205(.A1(new_n617), .A2(new_n621), .A3(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT83), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n617), .A2(new_n621), .A3(new_n633), .A4(new_n629), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n471), .A2(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  MUX2_X1   g219(.A(G99), .B(G111), .S(G2105), .Z(new_n645));
  AOI22_X1  g220(.A1(G123), .A2(new_n483), .B1(new_n645), .B2(G2104), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(new_n487), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT15), .B(G2435), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2427), .ZN(new_n655));
  INV_X1    g230(.A(G2430), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT84), .Z(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT17), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n669), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n671), .A3(new_n669), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n649), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n687), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G229));
  NOR2_X1   g277(.A1(G16), .A2(G19), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n569), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1341), .Z(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  OR2_X1    g282(.A1(G162), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(G35), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n708), .A2(KEYINPUT29), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(KEYINPUT29), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n706), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT100), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT23), .ZN(new_n716));
  INV_X1    g291(.A(G299), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n714), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1956), .Z(new_n719));
  INV_X1    g294(.A(KEYINPUT100), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(new_n706), .C1(new_n710), .C2(new_n711), .ZN(new_n721));
  AND4_X1   g296(.A1(new_n705), .A2(new_n713), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n471), .A2(G140), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  MUX2_X1   g299(.A(G104), .B(G116), .S(G2105), .Z(new_n725));
  AOI22_X1  g300(.A1(G128), .A2(new_n483), .B1(new_n725), .B2(G2104), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n707), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT93), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n707), .A2(G26), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT95), .B(G2067), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  AND2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  NOR2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n707), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n481), .B2(new_n707), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT97), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G2084), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(G2084), .ZN(new_n741));
  NAND2_X1  g316(.A1(G168), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n742), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n734), .A2(new_n740), .A3(new_n741), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G5), .A2(G16), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT99), .Z(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G301), .B2(new_n714), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G27), .A2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G164), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT31), .B(G11), .Z(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT30), .B(G28), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n759), .B1(new_n707), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n707), .A2(G32), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n471), .A2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n483), .A2(G129), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n473), .A2(G105), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n761), .B1(new_n707), .B2(new_n648), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n754), .A2(new_n758), .A3(new_n772), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n710), .A2(new_n711), .A3(new_n706), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n473), .A2(new_n775), .A3(G103), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(KEYINPUT25), .ZN(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n776), .B(new_n778), .C1(new_n487), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g356(.A1(G115), .A2(G2104), .ZN(new_n782));
  INV_X1    g357(.A(G127), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n465), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n781), .B1(G2105), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G29), .B2(G33), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G2072), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G2072), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(new_n753), .B2(new_n752), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n746), .A2(new_n747), .ZN(new_n791));
  AND4_X1   g366(.A1(new_n773), .A2(new_n774), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT90), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n622), .B2(new_n714), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT91), .B(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n722), .A2(new_n749), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT34), .ZN(new_n799));
  NOR2_X1   g374(.A1(G6), .A2(G16), .ZN(new_n800));
  INV_X1    g375(.A(G305), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT32), .B(G1981), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G22), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G166), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1971), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n587), .A2(new_n590), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G16), .B2(G23), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT88), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT33), .B(G1976), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT89), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n812), .A2(new_n815), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n799), .B(new_n808), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G95), .B(G107), .S(G2105), .Z(new_n819));
  AOI22_X1  g394(.A1(G119), .A2(new_n483), .B1(new_n819), .B2(G2104), .ZN(new_n820));
  INV_X1    g395(.A(G131), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n487), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(G29), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT87), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT86), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n823), .B(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(G16), .A2(G24), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G290), .B2(new_n714), .ZN(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n818), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n812), .B(new_n815), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n799), .B1(new_n834), .B2(new_n808), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT36), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n808), .B1(new_n816), .B2(new_n817), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n818), .A4(new_n832), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n798), .B1(new_n836), .B2(new_n840), .ZN(G311));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n840), .ZN(new_n842));
  INV_X1    g417(.A(new_n798), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT101), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n845), .B(new_n798), .C1(new_n836), .C2(new_n840), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(G150));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n537), .B2(new_n539), .ZN(new_n849));
  INV_X1    g424(.A(G93), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OAI22_X1  g426(.A1(new_n521), .A2(new_n850), .B1(new_n851), .B2(new_n508), .ZN(new_n852));
  OAI21_X1  g427(.A(G860), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n540), .A2(G55), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n558), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(G651), .A2(new_n858), .B1(new_n566), .B2(G93), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n859), .A3(KEYINPUT102), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n849), .B2(new_n852), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n568), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n568), .B1(new_n862), .B2(new_n860), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n569), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n568), .A2(new_n860), .A3(new_n862), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT38), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g445(.A(G559), .B(new_n623), .C1(new_n866), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n865), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n623), .A2(G559), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n871), .A2(new_n876), .A3(new_n880), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n871), .A2(new_n876), .ZN(new_n883));
  AOI21_X1  g458(.A(G860), .B1(new_n883), .B2(KEYINPUT39), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n882), .A2(KEYINPUT104), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT104), .B1(new_n882), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n854), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(new_n854), .C1(new_n885), .C2(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G145));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  MUX2_X1   g467(.A(G106), .B(G118), .S(G2105), .Z(new_n893));
  AOI22_X1  g468(.A1(G130), .A2(new_n483), .B1(new_n893), .B2(G2104), .ZN(new_n894));
  INV_X1    g469(.A(G142), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n487), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n640), .B(new_n896), .Z(new_n897));
  XOR2_X1   g472(.A(new_n822), .B(KEYINPUT108), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n724), .A2(new_n726), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G164), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n768), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G162), .B(new_n481), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n648), .B(KEYINPUT106), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n908), .B2(new_n912), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI211_X1 g491(.A(KEYINPUT109), .B(new_n911), .C1(new_n908), .C2(new_n912), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n892), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g495(.A1(G290), .A2(new_n591), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n809), .A2(new_n606), .A3(new_n605), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G303), .A2(G305), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n801), .A2(G166), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n921), .A2(new_n924), .A3(new_n922), .A4(new_n925), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n920), .B1(new_n929), .B2(KEYINPUT110), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(new_n931), .A3(new_n928), .A4(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n622), .A2(G299), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n617), .A2(new_n621), .A3(new_n717), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n872), .A2(new_n632), .A3(new_n634), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n872), .B1(new_n632), .B2(new_n634), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n872), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n635), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n934), .A2(new_n943), .A3(new_n935), .ZN(new_n944));
  INV_X1    g519(.A(new_n935), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n717), .B1(new_n617), .B2(new_n621), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT41), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n942), .A2(new_n937), .A3(new_n944), .A4(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n933), .A2(new_n940), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n940), .A2(new_n948), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n932), .A3(new_n930), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n933), .A2(new_n940), .A3(new_n948), .A4(KEYINPUT111), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G868), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n849), .A2(new_n852), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(G868), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT112), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n961), .B(new_n958), .C1(new_n955), .C2(G868), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n959), .ZN(G331));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n947), .A2(new_n944), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n540), .A2(G51), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n967), .A2(new_n535), .B1(new_n543), .B2(new_n547), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n531), .A2(new_n534), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n540), .A2(G51), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n544), .A3(new_n548), .A4(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n968), .B(new_n971), .C1(new_n863), .C2(new_n864), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n971), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n868), .A2(new_n973), .A3(new_n869), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n966), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n945), .A2(new_n946), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n972), .A3(new_n974), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n929), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n979), .A2(new_n892), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(KEYINPUT114), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n977), .A2(new_n972), .A3(new_n982), .A4(new_n974), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n947), .A2(KEYINPUT113), .A3(new_n944), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(new_n975), .C1(KEYINPUT113), .C2(new_n947), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n929), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n980), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT115), .B(new_n929), .C1(new_n984), .C2(new_n986), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n965), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  INV_X1    g567(.A(new_n929), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n947), .A2(new_n944), .B1(new_n972), .B2(new_n974), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n977), .A2(new_n972), .A3(new_n974), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n980), .A2(KEYINPUT43), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n989), .B2(new_n990), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n996), .A2(new_n979), .A3(new_n965), .A4(new_n892), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n992), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n998), .A2(new_n1005), .ZN(G397));
  NAND2_X1  g581(.A1(new_n501), .A2(new_n503), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT70), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n479), .B2(G114), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n492), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g586(.A1(G126), .A2(new_n483), .B1(new_n1011), .B2(new_n491), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n480), .A2(new_n468), .A3(G40), .A4(new_n474), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(G290), .B(G1986), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n900), .A2(G2067), .ZN(new_n1021));
  INV_X1    g596(.A(G2067), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n724), .A2(new_n1022), .A3(new_n726), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1996), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n768), .B(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n822), .A2(new_n825), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n822), .A2(new_n825), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1019), .B1(new_n1020), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  INV_X1    g607(.A(G1981), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n597), .A2(new_n601), .A3(new_n1033), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1035));
  INV_X1    g610(.A(G48), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1035), .A2(new_n508), .B1(new_n1036), .B2(new_n538), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n566), .A2(G86), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1034), .B1(new_n1039), .B2(KEYINPUT121), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  INV_X1    g616(.A(G86), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n601), .B1(new_n1042), .B2(new_n521), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1041), .B1(new_n1043), .B2(G1981), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1032), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(KEYINPUT121), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1041), .A3(G1981), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1032), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1034), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT119), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1052), .B(G1384), .C1(new_n1007), .C2(new_n1012), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1018), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1045), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n809), .A2(G1976), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n592), .A2(new_n1062), .A3(new_n594), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1056), .A2(new_n1061), .A3(new_n1063), .A4(new_n1058), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1018), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1384), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1971), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(KEYINPUT118), .A3(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1018), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1052), .B1(G164), .B2(G1384), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1070), .A2(KEYINPUT119), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1081), .A2(KEYINPUT120), .A3(new_n1083), .A4(new_n1082), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n706), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1050), .B1(new_n1078), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G303), .A2(G8), .ZN(new_n1091));
  XOR2_X1   g666(.A(new_n1091), .B(KEYINPUT55), .Z(new_n1092));
  AOI21_X1  g667(.A(new_n1065), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  INV_X1    g669(.A(G2084), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT120), .B1(new_n1054), .B2(new_n1082), .ZN(new_n1096));
  NOR4_X1   g671(.A1(new_n1051), .A2(new_n1053), .A3(new_n1085), .A4(KEYINPUT50), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1095), .B(new_n1079), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1054), .A2(KEYINPUT45), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1055), .A2(new_n1067), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n747), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1050), .B(G286), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1091), .B(KEYINPUT55), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1081), .A2(KEYINPUT50), .A3(new_n1083), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1015), .A2(new_n1082), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1018), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1106), .A2(new_n706), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1103), .B1(new_n1107), .B2(new_n1050), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1093), .A2(new_n1094), .A3(new_n1102), .A4(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1072), .A2(KEYINPUT118), .A3(new_n1073), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT118), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(G2090), .B(new_n1080), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1092), .B(G8), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1057), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1102), .A3(new_n1115), .A4(new_n1108), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT123), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1109), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(G8), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1120), .B2(new_n1103), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(new_n1093), .A3(new_n1102), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT124), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1121), .A2(new_n1093), .A3(new_n1124), .A4(new_n1102), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1119), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(G286), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1098), .A2(G168), .A3(new_n1101), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G8), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1130), .B2(G8), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(new_n1136), .C1(new_n1131), .C2(new_n1129), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1066), .A2(new_n1069), .A3(new_n757), .A4(new_n1071), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1100), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1139), .A2(G2078), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1141), .B(new_n1142), .C1(new_n1054), .C2(KEYINPUT45), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1079), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n753), .ZN(new_n1147));
  AOI21_X1  g722(.A(G301), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AND4_X1   g723(.A1(new_n1114), .A2(new_n1148), .A3(new_n1115), .A4(new_n1108), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1134), .A2(new_n1137), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1114), .A2(new_n1065), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1057), .A2(new_n1062), .A3(new_n595), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1034), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1056), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT56), .B(G2072), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1066), .A2(new_n1069), .A3(new_n1071), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1106), .B2(G1956), .ZN(new_n1157));
  AND3_X1   g732(.A1(G299), .A2(KEYINPUT125), .A3(KEYINPUT57), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT125), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1160), .B(new_n1156), .C1(G1956), .C2(new_n1106), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1162), .A2(KEYINPUT61), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1081), .A2(new_n1055), .A3(new_n1083), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(G2067), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1088), .B2(G1348), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n622), .A2(KEYINPUT60), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1066), .A2(new_n1069), .A3(new_n1025), .A4(new_n1071), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1174), .B2(new_n569), .ZN(new_n1175));
  AOI211_X1 g750(.A(KEYINPUT59), .B(new_n568), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1168), .A2(new_n1169), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT61), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1164), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(G1348), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1166), .B1(new_n1146), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n622), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n622), .B(new_n1167), .C1(new_n1088), .C2(G1348), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT60), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1181), .B2(new_n622), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1168), .A2(KEYINPUT126), .A3(new_n623), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n1162), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1179), .A2(new_n1185), .B1(new_n1189), .B2(new_n1163), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1088), .A2(G1961), .ZN(new_n1191));
  OAI21_X1  g766(.A(G171), .B1(new_n1191), .B2(new_n1144), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n467), .A2(G2105), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(G40), .A3(new_n474), .A4(new_n1142), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1139), .A2(new_n1138), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1147), .A2(G301), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1192), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT127), .B(KEYINPUT54), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT54), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1197), .B1(new_n1088), .B2(G1961), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1201), .B1(new_n1202), .B2(G171), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1145), .A2(new_n1147), .A3(G301), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1199), .A2(new_n1200), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1114), .A2(new_n1115), .A3(new_n1108), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1135), .B1(new_n1131), .B2(new_n1129), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1150), .B(new_n1154), .C1(new_n1190), .C2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1030), .B1(new_n1126), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(G290), .A2(G1986), .ZN(new_n1211));
  AOI21_X1  g786(.A(KEYINPUT48), .B1(new_n1211), .B2(new_n1019), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1211), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT48), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1019), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI211_X1 g791(.A(new_n1212), .B(new_n1216), .C1(new_n1019), .C2(new_n1029), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1024), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1019), .B1(new_n1218), .B2(new_n768), .ZN(new_n1219));
  NOR3_X1   g794(.A1(new_n1215), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT46), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1221), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1219), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g798(.A(new_n1223), .B(KEYINPUT47), .Z(new_n1224));
  NAND2_X1  g799(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1023), .B1(new_n1225), .B2(new_n1027), .ZN(new_n1226));
  AOI211_X1 g801(.A(new_n1217), .B(new_n1224), .C1(new_n1019), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1210), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g803(.A1(G401), .A2(G227), .A3(new_n460), .A4(G229), .ZN(new_n1230));
  NAND4_X1  g804(.A1(new_n991), .A2(new_n918), .A3(new_n997), .A4(new_n1230), .ZN(G225));
  INV_X1    g805(.A(G225), .ZN(G308));
endmodule


