//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT65), .B1(new_n207), .B2(G134gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n210));
  XNOR2_X1  g009(.A(G127gat), .B(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n211), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n213), .B(new_n208), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n216), .B(new_n219), .C1(new_n220), .C2(KEYINPUT2), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT70), .B(G141gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n217), .A3(new_n218), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n228), .A2(new_n216), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n221), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n215), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(KEYINPUT4), .B2(new_n231), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT70), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G141gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(G148gat), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n240), .A2(new_n223), .B1(new_n216), .B2(new_n228), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n216), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(G148gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n244), .B2(new_n227), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT3), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n221), .B(new_n247), .C1(new_n226), .C2(new_n229), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n215), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n235), .A2(KEYINPUT5), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n233), .B1(new_n215), .B2(new_n230), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n241), .A2(new_n245), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n212), .A4(new_n214), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT72), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(new_n233), .C1(new_n215), .C2(new_n230), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(new_n250), .A3(new_n249), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n254), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n249), .A2(new_n250), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n258), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT73), .A4(new_n261), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n215), .B(new_n230), .ZN(new_n268));
  INV_X1    g067(.A(new_n250), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n206), .B(new_n253), .C1(new_n267), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n206), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n263), .B2(new_n266), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n252), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT6), .B(new_n273), .C1(new_n274), .C2(new_n252), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G211gat), .A2(G218gat), .ZN(new_n280));
  INV_X1    g079(.A(G211gat), .ZN(new_n281));
  INV_X1    g080(.A(G218gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(G197gat), .A2(G204gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G197gat), .A2(G204gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n280), .B(new_n283), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n280), .ZN(new_n289));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(new_n287), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(KEYINPUT24), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT24), .A3(new_n296), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT25), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n298), .ZN(new_n308));
  AND2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n309), .A2(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  AND4_X1   g110(.A1(KEYINPUT25), .A2(new_n308), .A3(new_n306), .A4(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT27), .B1(new_n303), .B2(KEYINPUT64), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G183gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n304), .C1(KEYINPUT64), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(G190gat), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n316), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n299), .A2(KEYINPUT26), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n296), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n295), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(new_n299), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n307), .A2(new_n312), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT68), .B(KEYINPUT29), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n294), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n317), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n322), .A2(new_n325), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n308), .A2(new_n311), .A3(new_n306), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n306), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n329), .B(new_n293), .C1(new_n344), .C2(new_n328), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT69), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n350), .A3(new_n345), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT30), .A3(new_n353), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n346), .A2(KEYINPUT30), .A3(new_n351), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n279), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359));
  INV_X1    g158(.A(G50gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT76), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT75), .B(KEYINPUT31), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT77), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT82), .B(G22gat), .Z(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n288), .B2(new_n292), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n247), .B1(new_n367), .B2(KEYINPUT80), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  AOI211_X1 g168(.A(new_n369), .B(KEYINPUT29), .C1(new_n288), .C2(new_n292), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n230), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n293), .B1(new_n248), .B2(new_n331), .ZN(new_n372));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n374), .A3(KEYINPUT81), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n373), .B(KEYINPUT78), .Z(new_n380));
  INV_X1    g179(.A(new_n292), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n289), .B1(new_n291), .B2(new_n290), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n331), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT3), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n293), .A2(KEYINPUT79), .A3(new_n331), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n256), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n387), .B2(new_n372), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n366), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n371), .A2(KEYINPUT81), .A3(new_n374), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT81), .B1(new_n371), .B2(new_n374), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n388), .B(new_n366), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n365), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G22gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n392), .A3(new_n364), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n327), .A2(new_n215), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n338), .A2(new_n343), .A3(new_n212), .A4(new_n214), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G227gat), .ZN(new_n402));
  INV_X1    g201(.A(G233gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT66), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT66), .ZN(new_n406));
  INV_X1    g205(.A(new_n404), .ZN(new_n407));
  AOI211_X1 g206(.A(new_n406), .B(new_n407), .C1(new_n399), .C2(new_n400), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT32), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n405), .B2(new_n408), .ZN(new_n411));
  XOR2_X1   g210(.A(G15gat), .B(G43gat), .Z(new_n412));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT67), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(new_n401), .B2(new_n404), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT34), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n414), .ZN(new_n420));
  OAI221_X1 g219(.A(KEYINPUT32), .B1(new_n410), .B2(new_n420), .C1(new_n405), .C2(new_n408), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n415), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n415), .B2(new_n421), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n398), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT35), .B1(new_n358), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT88), .B(KEYINPUT35), .C1(new_n358), .C2(new_n424), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n356), .B1(new_n277), .B2(new_n278), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n415), .A2(new_n421), .ZN(new_n430));
  INV_X1    g229(.A(new_n419), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n419), .A3(new_n421), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT35), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n429), .A2(new_n434), .A3(new_n435), .A4(new_n398), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT87), .ZN(new_n437));
  INV_X1    g236(.A(new_n424), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n435), .A4(new_n429), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n427), .A2(new_n428), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT40), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n234), .B(new_n249), .C1(KEYINPUT4), .C2(new_n231), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n269), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n206), .B1(new_n445), .B2(KEYINPUT39), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT39), .B1(new_n268), .B2(new_n269), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n269), .B2(new_n444), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n442), .A2(KEYINPUT40), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n275), .A3(new_n356), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n453));
  NAND3_X1  g252(.A1(new_n333), .A2(new_n345), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n454), .B(KEYINPUT86), .Z(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n293), .B1(new_n330), .B2(new_n332), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n329), .B(new_n294), .C1(new_n344), .C2(new_n328), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(KEYINPUT37), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT84), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n455), .A2(new_n456), .A3(new_n351), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n350), .B1(new_n346), .B2(KEYINPUT37), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n353), .B(new_n461), .C1(new_n463), .C2(new_n456), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n398), .B(new_n452), .C1(new_n464), .C2(new_n279), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n434), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n432), .A2(KEYINPUT36), .A3(new_n433), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n366), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n395), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n392), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n392), .A2(new_n364), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n473), .A2(new_n365), .B1(new_n474), .B2(new_n396), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n358), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n441), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n479));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n481));
  NAND2_X1  g280(.A1(G29gat), .A2(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT90), .B(KEYINPUT15), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n480), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n494), .A3(new_n487), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(new_n482), .ZN(new_n496));
  OAI221_X1 g295(.A(KEYINPUT17), .B1(new_n483), .B2(new_n491), .C1(new_n496), .C2(new_n481), .ZN(new_n497));
  INV_X1    g296(.A(G22gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G15gat), .ZN(new_n499));
  INV_X1    g298(.A(G15gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G22gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G1gat), .ZN(new_n503));
  OR2_X1    g302(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(KEYINPUT16), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND4_X1   g309(.A1(new_n507), .A2(new_n509), .A3(new_n499), .A4(new_n501), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT93), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n506), .B(new_n514), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n483), .A2(new_n491), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n481), .B1(new_n495), .B2(new_n482), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n509), .A2(new_n499), .A3(new_n501), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n508), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G8gat), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n497), .A2(new_n516), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n515), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n507), .A3(new_n509), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n514), .B1(new_n528), .B2(new_n506), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n518), .A2(new_n519), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n524), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n479), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G197gat), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT11), .B(G169gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT12), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n535), .A2(new_n536), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n524), .A2(new_n533), .A3(KEYINPUT18), .A4(new_n534), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n516), .A2(new_n531), .A3(new_n523), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n533), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n534), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n535), .A2(new_n536), .B1(new_n547), .B2(new_n548), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(new_n545), .C1(new_n537), .C2(new_n542), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G120gat), .B(G148gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(G176gat), .B(G204gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT104), .Z(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n560), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT99), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n568), .A2(new_n570), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT100), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(G57gat), .A2(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G57gat), .A2(G64gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n589), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n587), .B(new_n596), .C1(new_n599), .C2(KEYINPUT96), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT10), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n574), .A2(new_n569), .A3(new_n575), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n582), .B1(KEYINPUT101), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n568), .A2(KEYINPUT101), .A3(new_n570), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n601), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n593), .A2(new_n600), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n578), .A2(new_n609), .A3(new_n581), .A4(new_n583), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT102), .B(KEYINPUT10), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n603), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT105), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n612), .B1(new_n608), .B2(new_n610), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n618), .B(new_n615), .C1(new_n619), .C2(new_n603), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n611), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n616), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n558), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n557), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g426(.A1(new_n609), .A2(new_n578), .A3(new_n581), .A4(new_n583), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n604), .A2(KEYINPUT101), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n579), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n609), .B1(new_n630), .B2(new_n606), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n613), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n603), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(KEYINPUT103), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n619), .B2(new_n603), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n636), .A3(new_n615), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n627), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n625), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n516), .A2(new_n523), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n645), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n657));
  XOR2_X1   g456(.A(G134gat), .B(G162gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n497), .A2(new_n520), .A3(new_n584), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G190gat), .B(G218gat), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n584), .B2(new_n531), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  INV_X1    g466(.A(new_n665), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(new_n661), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n660), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n663), .B1(new_n662), .B2(new_n665), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n667), .A3(new_n661), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n659), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n554), .A2(new_n639), .A3(new_n653), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n478), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n279), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n503), .ZN(G1324gat));
  INV_X1    g479(.A(G8gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n676), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n356), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT16), .B(G8gat), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n676), .A2(new_n357), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT42), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(KEYINPUT42), .B2(new_n685), .ZN(G1325gat));
  AOI21_X1  g486(.A(G15gat), .B1(new_n682), .B2(new_n434), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n469), .A2(G15gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT107), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n682), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n398), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n670), .A2(new_n673), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n441), .B2(new_n477), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n554), .A2(new_n639), .A3(new_n652), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n678), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n485), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT44), .B1(new_n478), .B2(new_n674), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  AOI211_X1 g502(.A(new_n703), .B(new_n695), .C1(new_n441), .C2(new_n477), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n705), .A2(new_n699), .A3(new_n697), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n701), .B1(new_n485), .B2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n698), .A2(new_n486), .A3(new_n356), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n705), .A2(new_n356), .A3(new_n697), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n486), .B2(new_n711), .ZN(G1329gat));
  NAND2_X1  g511(.A1(new_n478), .A2(new_n674), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n703), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n469), .A3(new_n715), .A4(new_n697), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n698), .A2(new_n719), .A3(new_n434), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  NAND4_X1  g522(.A1(new_n714), .A2(new_n475), .A3(new_n715), .A4(new_n697), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G50gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT48), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n698), .A2(new_n360), .A3(new_n475), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(new_n728), .C1(new_n726), .C2(KEYINPUT48), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n653), .A2(new_n674), .ZN(new_n733));
  AND4_X1   g532(.A1(new_n478), .A2(new_n554), .A3(new_n733), .A4(new_n639), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n699), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n356), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g539(.A(new_n434), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n434), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(G71gat), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n469), .A2(G71gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n734), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n475), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  INV_X1    g551(.A(new_n554), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n652), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n478), .A2(new_n674), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n754), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n696), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n678), .A2(G85gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n760), .A2(new_n639), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n639), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n753), .A2(new_n652), .A3(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n705), .A2(new_n699), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n766), .B2(new_n564), .ZN(G1336gat));
  NAND4_X1  g566(.A1(new_n714), .A2(new_n356), .A3(new_n715), .A4(new_n765), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n705), .A2(KEYINPUT114), .A3(new_n356), .A4(new_n765), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n356), .A2(new_n639), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n761), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n757), .A2(KEYINPUT113), .A3(new_n759), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n755), .A2(new_n779), .A3(new_n756), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n768), .A2(G92gat), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n783), .ZN(G1337gat));
  NOR2_X1   g583(.A1(new_n741), .A2(G99gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n760), .A2(new_n639), .A3(new_n761), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n714), .A2(new_n469), .A3(new_n715), .A4(new_n765), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G99gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(KEYINPUT115), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1338gat));
  NOR2_X1   g592(.A1(new_n398), .A2(G106gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n639), .A3(new_n780), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n714), .A2(new_n475), .A3(new_n715), .A4(new_n765), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n760), .A2(new_n639), .A3(new_n761), .A4(new_n794), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n797), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(G1339gat));
  AND3_X1   g602(.A1(new_n733), .A2(new_n554), .A3(new_n764), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n547), .A2(new_n548), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n534), .B1(new_n524), .B2(new_n533), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n541), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n552), .A2(new_n542), .A3(new_n545), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n639), .A2(new_n695), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n632), .A2(new_n633), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n618), .B1(new_n811), .B2(new_n615), .ZN(new_n812));
  INV_X1    g611(.A(new_n620), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n810), .B1(new_n614), .B2(new_n616), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n637), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n626), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n551), .A2(new_n553), .A3(new_n695), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n808), .A2(new_n807), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n674), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n819), .A2(new_n638), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n818), .B1(new_n637), .B2(new_n815), .ZN(new_n824));
  AND4_X1   g623(.A1(KEYINPUT116), .A2(new_n824), .A3(new_n814), .A4(new_n626), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n557), .B1(new_n621), .B2(new_n810), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT116), .B1(new_n826), .B2(new_n824), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n809), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n804), .B1(new_n829), .B2(new_n653), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n830), .A2(new_n356), .A3(new_n424), .A4(new_n678), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n753), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n639), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n652), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g636(.A(new_n695), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n839), .B(new_n840), .Z(G1343gat));
  NOR2_X1   g640(.A1(new_n830), .A2(new_n398), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n678), .A2(new_n469), .A3(new_n356), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n843), .A2(new_n845), .A3(G141gat), .A4(new_n554), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(KEYINPUT58), .ZN(new_n847));
  INV_X1    g646(.A(new_n225), .ZN(new_n848));
  XOR2_X1   g647(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n830), .B2(new_n398), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n826), .A2(new_n824), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n826), .A2(KEYINPUT116), .A3(new_n824), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n820), .A2(new_n822), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n817), .A2(new_n818), .B1(new_n637), .B2(new_n627), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n652), .B1(new_n860), .B2(new_n809), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n852), .B(new_n475), .C1(new_n861), .C2(new_n804), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n862), .A3(new_n844), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n848), .B1(new_n863), .B2(new_n554), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n862), .A3(KEYINPUT118), .A4(new_n844), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n753), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n846), .B1(new_n869), .B2(new_n848), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n865), .B(KEYINPUT119), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1344gat));
  NOR2_X1   g675(.A1(new_n843), .A2(new_n845), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n222), .A3(new_n639), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n844), .A2(new_n639), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n843), .A2(new_n852), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n842), .A2(new_n850), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n222), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n867), .A2(new_n639), .A3(new_n868), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(new_n879), .A3(G148gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n878), .B1(new_n887), .B2(new_n889), .ZN(G1345gat));
  NAND3_X1  g689(.A1(new_n877), .A2(new_n217), .A3(new_n652), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n867), .A2(new_n652), .A3(new_n868), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n217), .ZN(G1346gat));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n218), .A3(new_n674), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n867), .A2(new_n674), .A3(new_n868), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n218), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n357), .A2(new_n475), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n678), .A2(new_n742), .A3(new_n744), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n830), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(G169gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(new_n554), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n830), .A2(KEYINPUT121), .A3(new_n699), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT121), .B1(new_n830), .B2(new_n699), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n357), .B(new_n424), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n753), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n906), .B2(new_n901), .ZN(G1348gat));
  AOI21_X1  g706(.A(new_n424), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n774), .A2(G176gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G176gat), .B1(new_n900), .B2(new_n764), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1349gat));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n318), .A3(new_n652), .ZN(new_n913));
  OAI21_X1  g712(.A(G183gat), .B1(new_n900), .B2(new_n653), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g715(.A(new_n304), .B1(new_n899), .B2(new_n674), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n917), .A2(KEYINPUT123), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT124), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT123), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n917), .A2(new_n923), .A3(new_n918), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n919), .A2(new_n921), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n695), .A2(G190gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n905), .B2(new_n927), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n926), .A2(new_n908), .A3(new_n356), .A4(new_n927), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n925), .B(new_n932), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1351gat));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n470), .A2(new_n356), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n699), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT126), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n881), .A2(new_n882), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n935), .B1(new_n941), .B2(new_n554), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n882), .B2(new_n881), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(KEYINPUT127), .A3(new_n753), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n944), .A3(G197gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n903), .A2(new_n904), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n936), .A2(new_n398), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n554), .A2(G197gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  OR3_X1    g749(.A1(new_n948), .A2(G204gat), .A3(new_n764), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n941), .B2(new_n764), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  INV_X1    g754(.A(new_n948), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(new_n281), .A3(new_n652), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n943), .A2(new_n652), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n960));
  AOI211_X1 g759(.A(new_n960), .B(new_n281), .C1(new_n943), .C2(new_n652), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n959), .B2(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n941), .B2(new_n695), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n956), .A2(new_n282), .A3(new_n674), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


