

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XNOR2_X1 U323 ( .A(n330), .B(n329), .ZN(n344) );
  XNOR2_X1 U324 ( .A(n344), .B(n343), .ZN(n351) );
  XNOR2_X1 U325 ( .A(n420), .B(KEYINPUT48), .ZN(n559) );
  XNOR2_X1 U326 ( .A(n570), .B(KEYINPUT80), .ZN(n554) );
  AND2_X1 U327 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U328 ( .A(KEYINPUT74), .B(G64GAT), .Z(n292) );
  XOR2_X1 U329 ( .A(n333), .B(n384), .Z(n293) );
  NOR2_X1 U330 ( .A1(n409), .A2(n583), .ZN(n410) );
  AND2_X1 U331 ( .A1(n416), .A2(n415), .ZN(n417) );
  INV_X1 U332 ( .A(KEYINPUT122), .ZN(n435) );
  XNOR2_X1 U333 ( .A(n342), .B(n291), .ZN(n343) );
  NOR2_X1 U334 ( .A1(n481), .A2(n480), .ZN(n501) );
  NOR2_X1 U335 ( .A1(n478), .A2(n578), .ZN(n457) );
  NOR2_X1 U336 ( .A1(n561), .A2(n542), .ZN(n545) );
  XOR2_X1 U337 ( .A(n341), .B(n340), .Z(n519) );
  NOR2_X1 U338 ( .A1(n547), .A2(n458), .ZN(n463) );
  XOR2_X1 U339 ( .A(n432), .B(n431), .Z(n535) );
  XNOR2_X1 U340 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U341 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n295) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n310) );
  XOR2_X1 U345 ( .A(G176GAT), .B(KEYINPUT87), .Z(n297) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n303) );
  XOR2_X1 U348 ( .A(G183GAT), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U349 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n422) );
  XOR2_X1 U351 ( .A(n422), .B(KEYINPUT85), .Z(n301) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G71GAT), .Z(n392) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n304), .B(G127GAT), .ZN(n438) );
  XOR2_X1 U358 ( .A(n392), .B(n438), .Z(n306) );
  XNOR2_X1 U359 ( .A(G190GAT), .B(G134GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(n310), .B(n309), .Z(n538) );
  INV_X1 U363 ( .A(n538), .ZN(n547) );
  XOR2_X1 U364 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n312) );
  XNOR2_X1 U365 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U367 ( .A(KEYINPUT2), .B(n313), .Z(n442) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n342) );
  XNOR2_X1 U369 ( .A(G78GAT), .B(KEYINPUT70), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n314), .B(G148GAT), .ZN(n404) );
  XOR2_X1 U371 ( .A(n342), .B(n404), .Z(n316) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n442), .B(n317), .ZN(n328) );
  XOR2_X1 U375 ( .A(G204GAT), .B(KEYINPUT22), .Z(n319) );
  XNOR2_X1 U376 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U378 ( .A(n320), .B(G106GAT), .Z(n322) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G22GAT), .Z(n339) );
  XNOR2_X1 U380 ( .A(n339), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U382 ( .A(n323), .B(KEYINPUT23), .Z(n326) );
  XNOR2_X1 U383 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n324), .B(G211GAT), .ZN(n421) );
  XNOR2_X1 U385 ( .A(n421), .B(KEYINPUT91), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n478) );
  XOR2_X1 U388 ( .A(G29GAT), .B(G43GAT), .Z(n330) );
  XNOR2_X1 U389 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n329) );
  XOR2_X1 U390 ( .A(n344), .B(KEYINPUT67), .Z(n332) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n384) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G50GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n293), .B(n334), .ZN(n338) );
  XOR2_X1 U396 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n336) );
  XNOR2_X1 U397 ( .A(G113GAT), .B(G197GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U399 ( .A(n338), .B(n337), .Z(n341) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n428) );
  XNOR2_X1 U401 ( .A(n339), .B(n428), .ZN(n340) );
  XOR2_X1 U402 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n390) );
  XOR2_X1 U403 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n346) );
  XNOR2_X1 U404 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U406 ( .A(n347), .B(KEYINPUT10), .Z(n349) );
  XOR2_X1 U407 ( .A(G134GAT), .B(KEYINPUT78), .Z(n437) );
  XNOR2_X1 U408 ( .A(n437), .B(KEYINPUT79), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n365) );
  XOR2_X1 U411 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n363) );
  INV_X1 U412 ( .A(G99GAT), .ZN(n359) );
  INV_X1 U413 ( .A(KEYINPUT71), .ZN(n352) );
  NAND2_X1 U414 ( .A1(KEYINPUT72), .A2(n352), .ZN(n355) );
  INV_X1 U415 ( .A(KEYINPUT72), .ZN(n353) );
  NAND2_X1 U416 ( .A1(n353), .A2(KEYINPUT71), .ZN(n354) );
  NAND2_X1 U417 ( .A1(n355), .A2(n354), .ZN(n357) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G85GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n396) );
  XOR2_X1 U421 ( .A(G92GAT), .B(G218GAT), .Z(n361) );
  XNOR2_X1 U422 ( .A(G36GAT), .B(G190GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n424) );
  XNOR2_X1 U424 ( .A(n396), .B(n424), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n570) );
  NAND2_X1 U427 ( .A1(KEYINPUT36), .A2(n554), .ZN(n369) );
  INV_X1 U428 ( .A(KEYINPUT36), .ZN(n367) );
  INV_X1 U429 ( .A(n554), .ZN(n366) );
  NAND2_X1 U430 ( .A1(n367), .A2(n366), .ZN(n368) );
  NAND2_X1 U431 ( .A1(n369), .A2(n368), .ZN(n502) );
  XOR2_X1 U432 ( .A(G78GAT), .B(G211GAT), .Z(n371) );
  XNOR2_X1 U433 ( .A(G71GAT), .B(G155GAT), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U435 ( .A(G57GAT), .B(KEYINPUT13), .Z(n400) );
  XOR2_X1 U436 ( .A(n372), .B(n400), .Z(n374) );
  XNOR2_X1 U437 ( .A(G183GAT), .B(G127GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n388) );
  XOR2_X1 U439 ( .A(KEYINPUT14), .B(KEYINPUT84), .Z(n376) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n378) );
  XNOR2_X1 U443 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U445 ( .A(n380), .B(n379), .Z(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT82), .B(G64GAT), .Z(n382) );
  XNOR2_X1 U447 ( .A(G22GAT), .B(G8GAT), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(n388), .B(n387), .Z(n586) );
  NAND2_X1 U452 ( .A1(n502), .A2(n586), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n409) );
  XNOR2_X1 U454 ( .A(G176GAT), .B(G204GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n292), .B(n391), .ZN(n425) );
  XOR2_X1 U456 ( .A(n425), .B(n392), .Z(n394) );
  NAND2_X1 U457 ( .A1(G230GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U459 ( .A(n396), .B(n395), .Z(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n398) );
  XNOR2_X1 U461 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U463 ( .A(KEYINPUT32), .B(n399), .Z(n402) );
  XNOR2_X1 U464 ( .A(G92GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U466 ( .A(n403), .B(KEYINPUT69), .Z(n406) );
  XNOR2_X1 U467 ( .A(n404), .B(KEYINPUT68), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n583) );
  XNOR2_X1 U470 ( .A(KEYINPUT116), .B(n410), .ZN(n411) );
  AND2_X1 U471 ( .A1(n519), .A2(n411), .ZN(n412) );
  XNOR2_X1 U472 ( .A(KEYINPUT117), .B(n412), .ZN(n419) );
  INV_X1 U473 ( .A(n519), .ZN(n580) );
  XOR2_X1 U474 ( .A(n583), .B(KEYINPUT64), .Z(n413) );
  XNOR2_X1 U475 ( .A(n413), .B(KEYINPUT41), .ZN(n564) );
  NAND2_X1 U476 ( .A1(n580), .A2(n564), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n414), .B(KEYINPUT46), .ZN(n416) );
  NOR2_X1 U478 ( .A1(n570), .A2(n586), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n417), .B(KEYINPUT47), .ZN(n418) );
  NAND2_X1 U480 ( .A1(n419), .A2(n418), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U485 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U486 ( .A1(G226GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U488 ( .A(KEYINPUT121), .B(n535), .Z(n433) );
  NAND2_X1 U489 ( .A1(n559), .A2(n433), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n434), .B(KEYINPUT54), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n456) );
  XOR2_X1 U492 ( .A(G85GAT), .B(n437), .Z(n440) );
  XNOR2_X1 U493 ( .A(n438), .B(G162GAT), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n455) );
  XOR2_X1 U496 ( .A(G148GAT), .B(G120GAT), .Z(n444) );
  XNOR2_X1 U497 ( .A(G141GAT), .B(G29GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U502 ( .A(n448), .B(n447), .Z(n453) );
  XOR2_X1 U503 ( .A(KEYINPUT92), .B(G57GAT), .Z(n450) );
  NAND2_X1 U504 ( .A1(G225GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(n451), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U508 ( .A(n455), .B(n454), .Z(n532) );
  INV_X1 U509 ( .A(n532), .ZN(n487) );
  NAND2_X1 U510 ( .A1(n456), .A2(n487), .ZN(n578) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT55), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n463), .A2(n564), .ZN(n462) );
  XOR2_X1 U513 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n460) );
  XOR2_X1 U514 ( .A(G176GAT), .B(KEYINPUT56), .Z(n459) );
  XNOR2_X1 U515 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  NAND2_X1 U517 ( .A1(n463), .A2(n554), .ZN(n467) );
  XOR2_X1 U518 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n465) );
  INV_X1 U519 ( .A(G190GAT), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n489) );
  INV_X1 U521 ( .A(n535), .ZN(n491) );
  NOR2_X1 U522 ( .A1(n491), .A2(n547), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n478), .A2(n468), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT97), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT25), .ZN(n473) );
  NAND2_X1 U526 ( .A1(n547), .A2(n478), .ZN(n471) );
  XOR2_X1 U527 ( .A(n471), .B(KEYINPUT26), .Z(n558) );
  INV_X1 U528 ( .A(n558), .ZN(n579) );
  XOR2_X1 U529 ( .A(n535), .B(KEYINPUT27), .Z(n476) );
  NOR2_X1 U530 ( .A1(n579), .A2(n476), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n474), .A2(n532), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(n475), .ZN(n481) );
  NOR2_X1 U534 ( .A1(n476), .A2(n487), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT95), .ZN(n561) );
  XOR2_X1 U536 ( .A(n478), .B(KEYINPUT28), .Z(n498) );
  INV_X1 U537 ( .A(n498), .ZN(n542) );
  NAND2_X1 U538 ( .A1(n545), .A2(n547), .ZN(n479) );
  XOR2_X1 U539 ( .A(KEYINPUT96), .B(n479), .Z(n480) );
  INV_X1 U540 ( .A(n586), .ZN(n482) );
  NOR2_X1 U541 ( .A1(n482), .A2(n554), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  NOR2_X1 U543 ( .A1(n501), .A2(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT99), .B(n485), .ZN(n520) );
  OR2_X1 U545 ( .A1(n519), .A2(n583), .ZN(n505) );
  NOR2_X1 U546 ( .A1(n520), .A2(n505), .ZN(n486) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(n486), .Z(n497) );
  NOR2_X1 U548 ( .A1(n487), .A2(n497), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n491), .A2(n497), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT102), .B(n492), .Z(n493) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n493), .ZN(G1325GAT) );
  NOR2_X1 U554 ( .A1(n497), .A2(n547), .ZN(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  NOR2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(n499), .Z(n500) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  XOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .Z(n508) );
  NOR2_X1 U562 ( .A1(n586), .A2(n501), .ZN(n503) );
  NAND2_X1 U563 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT37), .B(n504), .Z(n531) );
  NOR2_X1 U565 ( .A1(n531), .A2(n505), .ZN(n506) );
  XNOR2_X2 U566 ( .A(n506), .B(KEYINPUT38), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n514), .A2(n532), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  XOR2_X1 U569 ( .A(G36GAT), .B(KEYINPUT105), .Z(n510) );
  NAND2_X1 U570 ( .A1(n514), .A2(n535), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1329GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n512) );
  NAND2_X1 U573 ( .A1(n538), .A2(n514), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U575 ( .A(n513), .B(G43GAT), .Z(G1330GAT) );
  XOR2_X1 U576 ( .A(G50GAT), .B(KEYINPUT107), .Z(n516) );
  NAND2_X1 U577 ( .A1(n514), .A2(n542), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n516), .B(n515), .ZN(G1331GAT) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n517), .B(KEYINPUT108), .ZN(n518) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(n518), .Z(n522) );
  NAND2_X1 U582 ( .A1(n564), .A2(n519), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n520), .A2(n530), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n527), .A2(n532), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U586 ( .A1(n535), .A2(n527), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT110), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G64GAT), .B(n524), .ZN(G1333GAT) );
  XOR2_X1 U589 ( .A(G71GAT), .B(KEYINPUT111), .Z(n526) );
  NAND2_X1 U590 ( .A1(n527), .A2(n538), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n542), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n534) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n541), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1336GAT) );
  XOR2_X1 U599 ( .A(G92GAT), .B(KEYINPUT113), .Z(n537) );
  NAND2_X1 U600 ( .A1(n541), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n541), .A2(n538), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT114), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G99GAT), .B(n540), .ZN(G1338GAT) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n543), .B(KEYINPUT44), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT118), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n559), .A2(n545), .ZN(n546) );
  NOR2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n580), .A2(n555), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U614 ( .A1(n555), .A2(n564), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U616 ( .A1(n555), .A2(n586), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT50), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  XOR2_X1 U622 ( .A(G141GAT), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n571), .A2(n580), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n566) );
  NAND2_X1 U628 ( .A1(n571), .A2(n564), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n567), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n571), .A2(n586), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT120), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G155GAT), .B(n569), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n463), .A2(n580), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n463), .A2(n586), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(n577), .Z(n582) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n589) );
  NAND2_X1 U645 ( .A1(n589), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U648 ( .A1(n589), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U651 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n502), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

