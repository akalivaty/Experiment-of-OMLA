//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT64), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(new_n468), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n477), .B(new_n480), .C1(G136), .C2(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT65), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT66), .A2(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n496), .B(new_n497), .C1(new_n485), .C2(new_n484), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n461), .A2(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n465), .B2(new_n466), .ZN(new_n500));
  INV_X1    g075(.A(new_n497), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT66), .A2(KEYINPUT4), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n498), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AND4_X1   g079(.A1(KEYINPUT67), .A2(new_n490), .A3(new_n494), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n493), .B1(new_n487), .B2(new_n489), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n506), .B2(new_n504), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(new_n513), .B1(G75), .B2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(KEYINPUT68), .A3(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n511), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(G543), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT69), .B(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n523), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n520), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n524), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n520), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n524), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT70), .Z(G188));
  AND2_X1   g131(.A1(new_n523), .A2(new_n511), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n534), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(G91), .A2(new_n557), .B1(new_n560), .B2(G651), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n562), .B(new_n563), .C1(new_n529), .C2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n564), .B1(KEYINPUT71), .B2(KEYINPUT9), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n520), .B(new_n566), .C1(KEYINPUT71), .C2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND2_X1  g148(.A1(new_n557), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n520), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  OAI21_X1  g152(.A(G61), .B1(new_n532), .B2(new_n533), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n578), .A2(new_n579), .B1(G73), .B2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n511), .A2(KEYINPUT73), .A3(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  AND2_X1   g158(.A1(KEYINPUT6), .A2(G651), .ZN(new_n584));
  NOR2_X1   g159(.A1(KEYINPUT6), .A2(G651), .ZN(new_n585));
  OAI211_X1 g160(.A(G48), .B(G543), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT74), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n520), .A2(new_n588), .A3(G48), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n587), .A2(new_n589), .B1(new_n557), .B2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n583), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n557), .A2(G85), .B1(G47), .B2(new_n520), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT75), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n510), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n523), .A2(new_n511), .A3(G92), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n534), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n568), .B(KEYINPUT72), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n550), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n604), .A2(new_n611), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT76), .ZN(G323));
  XOR2_X1   g191(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n617));
  XNOR2_X1  g192(.A(G323), .B(new_n617), .ZN(G282));
  NAND2_X1  g193(.A1(new_n467), .A2(new_n463), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n479), .A2(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n481), .B2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n622), .A2(G2100), .B1(new_n628), .B2(G2096), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G2100), .C2(new_n622), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT79), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT81), .Z(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n667), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n671), .C1(new_n664), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(new_n677), .Z(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  XNOR2_X1  g256(.A(KEYINPUT84), .B(G29), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G35), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G162), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT29), .B(G2090), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT25), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  AOI22_X1  g265(.A1(new_n481), .A2(G139), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n467), .A2(G127), .ZN(new_n693));
  NAND2_X1  g268(.A1(G115), .A2(G2104), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n461), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT92), .Z(new_n697));
  MUX2_X1   g272(.A(G33), .B(new_n697), .S(G29), .Z(new_n698));
  AOI21_X1  g273(.A(new_n686), .B1(G2072), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(G171), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G5), .B2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G28), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n705), .B2(KEYINPUT30), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(KEYINPUT30), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT31), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(G11), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G168), .A2(new_n700), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n700), .B2(G21), .ZN(new_n714));
  INV_X1    g289(.A(G1966), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n712), .B1(new_n628), .B2(new_n682), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n704), .B(new_n716), .C1(new_n715), .C2(new_n714), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n479), .A2(G129), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n463), .A2(G105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n481), .A2(G141), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n604), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G4), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n700), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n550), .B2(new_n700), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1341), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G34), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n740), .A2(new_n682), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G160), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n727), .ZN(new_n744));
  INV_X1    g319(.A(G2084), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n735), .A2(new_n738), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT91), .B(G2067), .Z(new_n748));
  AND2_X1   g323(.A1(new_n479), .A2(G128), .ZN(new_n749));
  NOR2_X1   g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT90), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n752));
  INV_X1    g327(.A(G140), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n468), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n682), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n748), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n756), .A2(new_n758), .A3(new_n748), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n759), .B(new_n760), .C1(new_n734), .C2(new_n733), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n699), .A2(new_n718), .A3(new_n747), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n702), .A2(new_n703), .B1(new_n745), .B2(new_n744), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n729), .B2(new_n730), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT97), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  NOR2_X1   g343(.A1(G164), .A2(new_n682), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G27), .B2(new_n682), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n763), .B(new_n767), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n698), .A2(G2072), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n700), .A2(G20), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT23), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n608), .B2(new_n700), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT98), .B(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n770), .A2(new_n768), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n778), .B(new_n779), .C1(new_n766), .C2(new_n765), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n762), .A2(new_n771), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G6), .B(G305), .S(G16), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT86), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT32), .B(G1981), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n700), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(G288), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n700), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n700), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n700), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT87), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n785), .B2(new_n784), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n792), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  MUX2_X1   g378(.A(G24), .B(G290), .S(G16), .Z(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(G1986), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(G1986), .ZN(new_n806));
  INV_X1    g381(.A(new_n682), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(G25), .ZN(new_n808));
  INV_X1    g383(.A(G131), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n461), .A2(G107), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n468), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n479), .B2(G119), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(new_n807), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT35), .B(G1991), .Z(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  NOR3_X1   g391(.A1(new_n805), .A2(new_n806), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n802), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(KEYINPUT36), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(KEYINPUT36), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT88), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n782), .B1(new_n820), .B2(new_n822), .ZN(G311));
  INV_X1    g398(.A(KEYINPUT89), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT88), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n821), .B(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n781), .B1(new_n825), .B2(new_n827), .ZN(G150));
  NAND2_X1  g403(.A1(new_n520), .A2(G55), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n524), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n510), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT101), .B(G860), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  INV_X1    g414(.A(new_n550), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n550), .B1(new_n833), .B2(new_n831), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n841), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n604), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n837), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n839), .B1(new_n852), .B2(new_n854), .ZN(G145));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n498), .B(new_n856), .C1(new_n500), .C2(new_n503), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n496), .B1(new_n484), .B2(new_n485), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT66), .B(KEYINPUT4), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n856), .B1(new_n861), .B2(new_n498), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n506), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g440(.A(KEYINPUT103), .B(new_n506), .C1(new_n858), .C2(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n749), .A2(new_n754), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n870), .A2(new_n871), .B1(new_n719), .B2(new_n725), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n755), .A2(new_n865), .A3(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n726), .A3(new_n869), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n872), .A2(new_n697), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n696), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n461), .B2(G118), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n878), .A2(new_n461), .A3(G118), .ZN(new_n881));
  INV_X1    g456(.A(G142), .ZN(new_n882));
  OAI22_X1  g457(.A1(new_n880), .A2(new_n881), .B1(new_n468), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n479), .B2(G130), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n620), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n813), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n875), .A2(new_n877), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n628), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G162), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n875), .B2(new_n877), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT105), .A4(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n889), .B1(new_n887), .B2(new_n890), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n895), .B2(new_n898), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT106), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT40), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n903), .A2(new_n906), .ZN(G395));
  XNOR2_X1  g482(.A(new_n846), .B(new_n614), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n608), .A2(new_n603), .ZN(new_n909));
  NOR2_X1   g484(.A1(G299), .A2(new_n604), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n909), .B2(new_n910), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n916), .B2(new_n908), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(G166), .B(KEYINPUT107), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G305), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n788), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n918), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G868), .B2(new_n836), .ZN(G295));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n836), .ZN(G331));
  XNOR2_X1  g502(.A(G286), .B(G171), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n846), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n841), .A3(new_n844), .A4(new_n845), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT108), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n847), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n916), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n931), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(new_n911), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n922), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n938), .B2(KEYINPUT109), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(new_n922), .A3(new_n940), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n937), .ZN(new_n942));
  INV_X1    g517(.A(new_n922), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n932), .A2(new_n934), .A3(new_n911), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n916), .A2(new_n936), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n941), .A4(new_n939), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n946), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n941), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n947), .A2(new_n948), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n947), .A2(new_n948), .B1(new_n916), .B2(new_n936), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n922), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n960), .C2(new_n963), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n957), .B1(new_n969), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n865), .A2(new_n971), .A3(new_n866), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT112), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n865), .A2(new_n975), .A3(new_n971), .A4(new_n866), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n470), .A2(new_n473), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n726), .B(G1996), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n868), .B(G2067), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n813), .A2(new_n815), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n813), .A2(new_n815), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(G290), .B(G1986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g565(.A1(G286), .A2(G8), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT119), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n504), .A2(KEYINPUT102), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n857), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n994), .B2(new_n506), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n980), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n490), .A2(new_n504), .A3(new_n494), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT67), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n506), .A2(KEYINPUT67), .A3(new_n504), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n971), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n997), .A2(new_n745), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n863), .A2(new_n971), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n980), .B1(new_n1005), .B2(new_n974), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n971), .A4(new_n1001), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1966), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n992), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(new_n979), .C1(KEYINPUT45), .C2(new_n995), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n715), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n997), .A2(new_n745), .A3(new_n1003), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1009), .B(KEYINPUT51), .C1(new_n1014), .C2(new_n992), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(new_n992), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1016), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n990), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n992), .B1(new_n1025), .B2(G8), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1020), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT120), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(KEYINPUT62), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n980), .B1(new_n1002), .B2(new_n974), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n865), .A2(KEYINPUT45), .A3(new_n971), .A4(new_n866), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n796), .ZN(new_n1034));
  INV_X1    g609(.A(G2090), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n997), .A2(new_n1035), .A3(new_n1003), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1010), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G166), .A2(new_n1010), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT55), .Z(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n589), .A2(new_n587), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n557), .A2(G86), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n510), .B1(new_n580), .B2(new_n581), .ZN(new_n1045));
  OAI21_X1  g620(.A(G1981), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1981), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n583), .A2(new_n590), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1048), .A3(KEYINPUT49), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n863), .A2(new_n979), .A3(new_n971), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(G8), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n788), .A2(G1976), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(G8), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1051), .A2(new_n1052), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1054), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n979), .B1(new_n995), .B2(new_n996), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1000), .A2(new_n996), .A3(new_n971), .A4(new_n1001), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n508), .A2(KEYINPUT114), .A3(new_n996), .A4(new_n971), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1035), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1010), .B1(new_n1070), .B2(new_n1034), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1041), .B(new_n1063), .C1(new_n1040), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1011), .B2(G2078), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1006), .A2(KEYINPUT121), .A3(new_n768), .A4(new_n1007), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(KEYINPUT53), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1031), .A2(new_n1032), .A3(new_n768), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n863), .A2(new_n996), .A3(new_n971), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n505), .A2(new_n507), .A3(G1384), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n979), .B(new_n1079), .C1(new_n1080), .C2(new_n996), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1077), .A2(new_n1078), .B1(new_n1081), .B2(new_n703), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1072), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1023), .A2(new_n1030), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1063), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1055), .B(new_n788), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1048), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(G8), .A3(new_n1050), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1017), .A2(G286), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1041), .A2(new_n1092), .A3(KEYINPUT63), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1036), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1971), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1039), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT115), .A3(new_n1063), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT115), .B1(new_n1097), .B2(new_n1063), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1092), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1072), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1091), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1086), .A2(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(new_n568), .B(KEYINPUT57), .Z(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1031), .A2(new_n1032), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1069), .B2(G1956), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1031), .A2(new_n1032), .A3(new_n1110), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1113), .A2(KEYINPUT116), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1068), .A2(new_n1067), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1064), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1113), .A2(KEYINPUT116), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n1107), .A3(new_n1121), .A4(new_n1111), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1115), .A2(new_n1122), .A3(KEYINPUT61), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1050), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1033), .A2(G1996), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT117), .A3(new_n550), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT59), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(KEYINPUT117), .A3(new_n1132), .A4(new_n550), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n603), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1050), .A2(G2067), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1081), .B2(new_n734), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT118), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1348), .B1(new_n997), .B2(new_n1003), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  NOR4_X1   g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1139), .A4(new_n1137), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1136), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n996), .B1(new_n508), .B2(new_n971), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1079), .A2(new_n979), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n734), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1137), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n1149), .A3(new_n1140), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1143), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1138), .A2(KEYINPUT118), .A3(new_n1140), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1136), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1145), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1125), .A2(new_n1126), .A3(new_n1134), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1115), .B1(new_n603), .B2(new_n1138), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1076), .A2(new_n1082), .A3(G301), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1076), .A2(new_n1082), .A3(KEYINPUT123), .A4(G301), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1162), .A2(KEYINPUT54), .A3(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1032), .A2(KEYINPUT53), .A3(new_n768), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n977), .A2(KEYINPUT122), .A3(new_n979), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT122), .B1(new_n977), .B2(new_n979), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1082), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(G171), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(G301), .A3(new_n1082), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1084), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1021), .A2(new_n1022), .A3(new_n1072), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1159), .A2(new_n1171), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n989), .B1(new_n1106), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n982), .A2(new_n983), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1179), .A2(new_n984), .B1(G2067), .B2(new_n755), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n981), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT124), .Z(new_n1182));
  OR2_X1    g757(.A1(new_n977), .A2(new_n980), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1183), .A2(G1986), .A3(G290), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT48), .Z(new_n1185));
  NAND2_X1  g760(.A1(new_n986), .A2(new_n981), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT126), .Z(new_n1187));
  AOI21_X1  g762(.A(new_n1182), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT46), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n983), .B(new_n726), .C1(new_n1189), .C2(G1996), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n981), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1189), .B1(new_n1183), .B2(G1996), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1192), .A2(KEYINPUT125), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1192), .A2(KEYINPUT125), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1191), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT47), .ZN(new_n1196));
  OR2_X1    g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1188), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT127), .B1(new_n1178), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1175), .A2(new_n1171), .A3(new_n1176), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1086), .A2(new_n1105), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n988), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1188), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1200), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g784(.A1(new_n946), .A2(new_n955), .ZN(new_n1211));
  OR2_X1    g785(.A1(G227), .A2(new_n459), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(G401), .A3(new_n1212), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n1211), .B(new_n1213), .C1(new_n900), .C2(new_n901), .ZN(G225));
  INV_X1    g788(.A(G225), .ZN(G308));
endmodule


