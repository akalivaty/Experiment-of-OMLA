

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U548 ( .A1(n740), .A2(G1996), .ZN(n718) );
  INV_X1 U549 ( .A(n761), .ZN(n740) );
  NAND2_X1 U550 ( .A1(n715), .A2(n714), .ZN(n761) );
  NOR2_X1 U551 ( .A1(G651), .A2(n614), .ZN(n639) );
  XNOR2_X1 U552 ( .A(G1341), .B(G2435), .ZN(n520) );
  XOR2_X1 U553 ( .A(G2451), .B(G2446), .Z(n512) );
  XNOR2_X1 U554 ( .A(G1348), .B(KEYINPUT101), .ZN(n511) );
  XNOR2_X1 U555 ( .A(n512), .B(n511), .ZN(n516) );
  XOR2_X1 U556 ( .A(G2430), .B(G2454), .Z(n514) );
  XNOR2_X1 U557 ( .A(G2427), .B(KEYINPUT100), .ZN(n513) );
  XNOR2_X1 U558 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U559 ( .A(n516), .B(n515), .Z(n518) );
  XNOR2_X1 U560 ( .A(G2443), .B(G2438), .ZN(n517) );
  XNOR2_X1 U561 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U562 ( .A(n520), .B(n519), .ZN(n521) );
  AND2_X1 U563 ( .A1(n521), .A2(G14), .ZN(G401) );
  AND2_X1 U564 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U565 ( .A(G57), .ZN(G237) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n522), .Z(n989) );
  NAND2_X1 U568 ( .A1(G137), .A2(n989), .ZN(n524) );
  INV_X1 U569 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n527), .ZN(n985) );
  NAND2_X1 U571 ( .A1(G125), .A2(n985), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n532) );
  NAND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U574 ( .A(n525), .B(KEYINPUT65), .ZN(n986) );
  NAND2_X1 U575 ( .A1(G113), .A2(n986), .ZN(n526) );
  XNOR2_X1 U576 ( .A(n526), .B(KEYINPUT66), .ZN(n530) );
  AND2_X1 U577 ( .A1(n527), .A2(G2104), .ZN(n990) );
  NAND2_X1 U578 ( .A1(G101), .A2(n990), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n679) );
  BUF_X1 U582 ( .A(n679), .Z(G160) );
  XNOR2_X1 U583 ( .A(KEYINPUT67), .B(G651), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G543), .A2(n535), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n533), .Z(n638) );
  NAND2_X1 U586 ( .A1(n638), .A2(G64), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT69), .ZN(n542) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U589 ( .A1(n633), .A2(G90), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n614) );
  NOR2_X1 U591 ( .A1(n614), .A2(n535), .ZN(n634) );
  NAND2_X1 U592 ( .A1(G77), .A2(n634), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n538), .B(KEYINPUT9), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G52), .A2(n639), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U597 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U598 ( .A1(G7), .A2(G661), .ZN(n543) );
  XNOR2_X1 U599 ( .A(n543), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U600 ( .A(G223), .ZN(n809) );
  NAND2_X1 U601 ( .A1(n809), .A2(G567), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT11), .B(n544), .Z(G234) );
  NAND2_X1 U603 ( .A1(n638), .A2(G56), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT14), .B(n545), .Z(n552) );
  NAND2_X1 U605 ( .A1(G81), .A2(n633), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n546), .B(KEYINPUT12), .ZN(n547) );
  XNOR2_X1 U607 ( .A(n547), .B(KEYINPUT72), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G68), .A2(n634), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT13), .B(n550), .Z(n551) );
  NOR2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n639), .A2(G43), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n949) );
  INV_X1 U614 ( .A(G860), .ZN(n588) );
  OR2_X1 U615 ( .A1(n949), .A2(n588), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT73), .B(n555), .Z(G153) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(G868), .A2(G301), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G54), .A2(n639), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G79), .A2(n634), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G66), .A2(n638), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n633), .A2(G92), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT74), .B(n558), .Z(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT15), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT75), .B(n564), .ZN(n823) );
  INV_X1 U629 ( .A(G868), .ZN(n653) );
  NAND2_X1 U630 ( .A1(n823), .A2(n653), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(G284) );
  NAND2_X1 U632 ( .A1(G89), .A2(n633), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT4), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT76), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G76), .A2(n634), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT5), .B(n571), .ZN(n577) );
  XNOR2_X1 U638 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n639), .A2(G51), .ZN(n573) );
  NAND2_X1 U640 ( .A1(G63), .A2(n638), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(n639), .A2(G53), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G65), .A2(n638), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n633), .A2(G91), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G78), .A2(n634), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n828) );
  INV_X1 U653 ( .A(n828), .ZN(G299) );
  NOR2_X1 U654 ( .A1(G286), .A2(n653), .ZN(n586) );
  NOR2_X1 U655 ( .A1(G868), .A2(G299), .ZN(n585) );
  NOR2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U657 ( .A(KEYINPUT78), .B(n587), .ZN(G297) );
  NAND2_X1 U658 ( .A1(n588), .A2(G559), .ZN(n589) );
  INV_X1 U659 ( .A(n823), .ZN(n946) );
  NAND2_X1 U660 ( .A1(n589), .A2(n946), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT16), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT79), .B(n591), .Z(G148) );
  NOR2_X1 U663 ( .A1(G868), .A2(n949), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G868), .A2(n946), .ZN(n592) );
  NOR2_X1 U665 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(G282) );
  XOR2_X1 U667 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n596) );
  NAND2_X1 U668 ( .A1(G123), .A2(n985), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U670 ( .A(n597), .B(KEYINPUT80), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n986), .A2(G111), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G135), .A2(n989), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G99), .A2(n990), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n974) );
  XNOR2_X1 U677 ( .A(G2096), .B(n974), .ZN(n605) );
  INV_X1 U678 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G559), .A2(n946), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n949), .B(n606), .ZN(n650) );
  NOR2_X1 U682 ( .A1(n650), .A2(G860), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n639), .A2(G55), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G67), .A2(n638), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n633), .A2(G93), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G80), .A2(n634), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n652) );
  XNOR2_X1 U690 ( .A(n613), .B(n652), .ZN(G145) );
  NAND2_X1 U691 ( .A1(G87), .A2(n614), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n638), .A2(n617), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n639), .A2(G49), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(G288) );
  NAND2_X1 U697 ( .A1(n633), .A2(G88), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G75), .A2(n634), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n639), .A2(G50), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G62), .A2(n638), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(G166) );
  NAND2_X1 U704 ( .A1(G86), .A2(n633), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G48), .A2(n639), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n634), .A2(G73), .ZN(n628) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n628), .Z(n629) );
  NOR2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G61), .A2(n638), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U712 ( .A1(n633), .A2(G85), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G72), .A2(n634), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT68), .B(n637), .Z(n643) );
  NAND2_X1 U716 ( .A1(n638), .A2(G60), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n639), .A2(G47), .ZN(n640) );
  AND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(G290) );
  XOR2_X1 U720 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n644) );
  XNOR2_X1 U721 ( .A(G288), .B(n644), .ZN(n645) );
  XOR2_X1 U722 ( .A(n645), .B(n652), .Z(n647) );
  XNOR2_X1 U723 ( .A(n828), .B(G166), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(G305), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n649), .B(G290), .ZN(n945) );
  XOR2_X1 U727 ( .A(n650), .B(n945), .Z(n651) );
  NAND2_X1 U728 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U731 ( .A(KEYINPUT83), .B(n656), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n657) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(KEYINPUT84), .B(G44), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n661), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U739 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  XNOR2_X1 U740 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U741 ( .A1(G219), .A2(G220), .ZN(n662) );
  XOR2_X1 U742 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U743 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U744 ( .A1(G96), .A2(n664), .ZN(n944) );
  NAND2_X1 U745 ( .A1(G2106), .A2(n944), .ZN(n665) );
  XNOR2_X1 U746 ( .A(KEYINPUT85), .B(n665), .ZN(n670) );
  NAND2_X1 U747 ( .A1(G120), .A2(G69), .ZN(n666) );
  NOR2_X1 U748 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U749 ( .A1(G108), .A2(n667), .ZN(n943) );
  NAND2_X1 U750 ( .A1(G567), .A2(n943), .ZN(n668) );
  XOR2_X1 U751 ( .A(KEYINPUT86), .B(n668), .Z(n669) );
  NOR2_X1 U752 ( .A1(n670), .A2(n669), .ZN(G319) );
  INV_X1 U753 ( .A(G319), .ZN(n1003) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n671) );
  NOR2_X1 U755 ( .A1(n1003), .A2(n671), .ZN(n814) );
  NAND2_X1 U756 ( .A1(n814), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(G138), .A2(n989), .ZN(n673) );
  NAND2_X1 U758 ( .A1(G102), .A2(n990), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G126), .A2(n985), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G114), .A2(n986), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U763 ( .A1(n677), .A2(n676), .ZN(G164) );
  XNOR2_X1 U764 ( .A(G166), .B(KEYINPUT87), .ZN(G303) );
  XNOR2_X1 U765 ( .A(G1986), .B(KEYINPUT88), .ZN(n678) );
  XNOR2_X1 U766 ( .A(n678), .B(G290), .ZN(n837) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n714) );
  NAND2_X1 U768 ( .A1(n679), .A2(G40), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n804) );
  NAND2_X1 U770 ( .A1(n837), .A2(n804), .ZN(n793) );
  NAND2_X1 U771 ( .A1(G140), .A2(n989), .ZN(n681) );
  NAND2_X1 U772 ( .A1(G104), .A2(n990), .ZN(n680) );
  NAND2_X1 U773 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n682), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT90), .B(KEYINPUT35), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n985), .A2(G128), .ZN(n685) );
  NAND2_X1 U777 ( .A1(n986), .A2(G116), .ZN(n683) );
  XOR2_X1 U778 ( .A(KEYINPUT89), .B(n683), .Z(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U780 ( .A(n687), .B(n686), .Z(n688) );
  NOR2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U782 ( .A(KEYINPUT36), .B(n690), .ZN(n982) );
  XNOR2_X1 U783 ( .A(G2067), .B(KEYINPUT37), .ZN(n802) );
  NOR2_X1 U784 ( .A1(n982), .A2(n802), .ZN(n691) );
  XOR2_X1 U785 ( .A(KEYINPUT91), .B(n691), .Z(n935) );
  NAND2_X1 U786 ( .A1(n804), .A2(n935), .ZN(n800) );
  NAND2_X1 U787 ( .A1(G129), .A2(n985), .ZN(n693) );
  NAND2_X1 U788 ( .A1(G117), .A2(n986), .ZN(n692) );
  NAND2_X1 U789 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n990), .A2(G105), .ZN(n694) );
  XOR2_X1 U791 ( .A(KEYINPUT38), .B(n694), .Z(n695) );
  NOR2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U793 ( .A(n697), .B(KEYINPUT94), .ZN(n699) );
  NAND2_X1 U794 ( .A1(G141), .A2(n989), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n980) );
  NAND2_X1 U796 ( .A1(n980), .A2(G1996), .ZN(n709) );
  NAND2_X1 U797 ( .A1(G131), .A2(n989), .ZN(n701) );
  NAND2_X1 U798 ( .A1(G95), .A2(n990), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U800 ( .A1(G119), .A2(n985), .ZN(n703) );
  NAND2_X1 U801 ( .A1(G107), .A2(n986), .ZN(n702) );
  NAND2_X1 U802 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U803 ( .A(KEYINPUT92), .B(n704), .ZN(n705) );
  NOR2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U805 ( .A(n707), .B(KEYINPUT93), .ZN(n976) );
  NAND2_X1 U806 ( .A1(n976), .A2(G1991), .ZN(n708) );
  AND2_X1 U807 ( .A1(n709), .A2(n708), .ZN(n929) );
  XNOR2_X1 U808 ( .A(KEYINPUT95), .B(n804), .ZN(n710) );
  NOR2_X1 U809 ( .A1(n929), .A2(n710), .ZN(n797) );
  INV_X1 U810 ( .A(n797), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n800), .A2(n711), .ZN(n791) );
  INV_X1 U812 ( .A(KEYINPUT96), .ZN(n712) );
  XNOR2_X1 U813 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U814 ( .A1(G8), .A2(n761), .ZN(n784) );
  NOR2_X1 U815 ( .A1(G1981), .A2(G305), .ZN(n716) );
  XOR2_X1 U816 ( .A(n716), .B(KEYINPUT24), .Z(n717) );
  NOR2_X1 U817 ( .A1(n784), .A2(n717), .ZN(n789) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n761), .ZN(n745) );
  NAND2_X1 U819 ( .A1(G8), .A2(n745), .ZN(n759) );
  NOR2_X1 U820 ( .A1(G1966), .A2(n784), .ZN(n757) );
  XOR2_X1 U821 ( .A(n718), .B(KEYINPUT26), .Z(n720) );
  NAND2_X1 U822 ( .A1(n761), .A2(G1341), .ZN(n719) );
  NAND2_X1 U823 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U824 ( .A1(n949), .A2(n721), .ZN(n725) );
  NAND2_X1 U825 ( .A1(G1348), .A2(n761), .ZN(n723) );
  NAND2_X1 U826 ( .A1(G2067), .A2(n740), .ZN(n722) );
  NAND2_X1 U827 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U828 ( .A1(n823), .A2(n726), .ZN(n724) );
  OR2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U830 ( .A1(n823), .A2(n726), .ZN(n727) );
  NAND2_X1 U831 ( .A1(n728), .A2(n727), .ZN(n733) );
  NAND2_X1 U832 ( .A1(n740), .A2(G2072), .ZN(n729) );
  XNOR2_X1 U833 ( .A(n729), .B(KEYINPUT27), .ZN(n731) );
  XNOR2_X1 U834 ( .A(G1956), .B(KEYINPUT97), .ZN(n858) );
  NOR2_X1 U835 ( .A1(n858), .A2(n740), .ZN(n730) );
  NOR2_X1 U836 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U837 ( .A1(n828), .A2(n734), .ZN(n732) );
  NAND2_X1 U838 ( .A1(n733), .A2(n732), .ZN(n737) );
  NOR2_X1 U839 ( .A1(n828), .A2(n734), .ZN(n735) );
  XOR2_X1 U840 ( .A(n735), .B(KEYINPUT28), .Z(n736) );
  NAND2_X1 U841 ( .A1(n737), .A2(n736), .ZN(n739) );
  XOR2_X1 U842 ( .A(KEYINPUT98), .B(KEYINPUT29), .Z(n738) );
  XNOR2_X1 U843 ( .A(n739), .B(n738), .ZN(n744) );
  XOR2_X1 U844 ( .A(G2078), .B(KEYINPUT25), .Z(n884) );
  NOR2_X1 U845 ( .A1(n884), .A2(n761), .ZN(n742) );
  NOR2_X1 U846 ( .A1(n740), .A2(G1961), .ZN(n741) );
  NOR2_X1 U847 ( .A1(n742), .A2(n741), .ZN(n750) );
  OR2_X1 U848 ( .A1(n750), .A2(G301), .ZN(n743) );
  NAND2_X1 U849 ( .A1(n744), .A2(n743), .ZN(n755) );
  NOR2_X1 U850 ( .A1(n757), .A2(n745), .ZN(n746) );
  NAND2_X1 U851 ( .A1(G8), .A2(n746), .ZN(n747) );
  XOR2_X1 U852 ( .A(KEYINPUT30), .B(n747), .Z(n749) );
  INV_X1 U853 ( .A(G168), .ZN(n748) );
  NAND2_X1 U854 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U855 ( .A1(n750), .A2(G301), .ZN(n751) );
  NAND2_X1 U856 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U857 ( .A(n753), .B(KEYINPUT31), .ZN(n754) );
  NAND2_X1 U858 ( .A1(n755), .A2(n754), .ZN(n760) );
  INV_X1 U859 ( .A(n760), .ZN(n756) );
  NOR2_X1 U860 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U861 ( .A1(n759), .A2(n758), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n760), .A2(G286), .ZN(n766) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n784), .ZN(n763) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U865 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U866 ( .A1(n764), .A2(G303), .ZN(n765) );
  NAND2_X1 U867 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U868 ( .A1(n767), .A2(G8), .ZN(n768) );
  XNOR2_X1 U869 ( .A(n768), .B(KEYINPUT32), .ZN(n769) );
  NAND2_X1 U870 ( .A1(n770), .A2(n769), .ZN(n783) );
  NOR2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n776) );
  NOR2_X1 U872 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U873 ( .A1(n776), .A2(n771), .ZN(n832) );
  NAND2_X1 U874 ( .A1(n783), .A2(n832), .ZN(n772) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n831) );
  NAND2_X1 U876 ( .A1(n772), .A2(n831), .ZN(n773) );
  NOR2_X1 U877 ( .A1(n784), .A2(n773), .ZN(n774) );
  XNOR2_X1 U878 ( .A(n774), .B(KEYINPUT64), .ZN(n775) );
  NOR2_X1 U879 ( .A1(KEYINPUT33), .A2(n775), .ZN(n779) );
  NAND2_X1 U880 ( .A1(n776), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U881 ( .A1(n777), .A2(n784), .ZN(n778) );
  NOR2_X1 U882 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U883 ( .A(G1981), .B(G305), .Z(n842) );
  NAND2_X1 U884 ( .A1(n780), .A2(n842), .ZN(n787) );
  NOR2_X1 U885 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U886 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U887 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U888 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U889 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U890 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U891 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n793), .A2(n792), .ZN(n807) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n980), .ZN(n923) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n795) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n976), .ZN(n794) );
  XOR2_X1 U896 ( .A(KEYINPUT99), .B(n794), .Z(n907) );
  NOR2_X1 U897 ( .A1(n795), .A2(n907), .ZN(n796) );
  NOR2_X1 U898 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U899 ( .A1(n923), .A2(n798), .ZN(n799) );
  XNOR2_X1 U900 ( .A(n799), .B(KEYINPUT39), .ZN(n801) );
  NAND2_X1 U901 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n982), .A2(n802), .ZN(n906) );
  NAND2_X1 U903 ( .A1(n803), .A2(n906), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n808), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n809), .ZN(G217) );
  INV_X1 U908 ( .A(G661), .ZN(n811) );
  NAND2_X1 U909 ( .A1(G2), .A2(G15), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U911 ( .A(KEYINPUT102), .B(n812), .Z(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n813) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(G188) );
  XNOR2_X1 U914 ( .A(G69), .B(KEYINPUT103), .ZN(G235) );
  NAND2_X1 U916 ( .A1(G136), .A2(n989), .ZN(n816) );
  NAND2_X1 U917 ( .A1(G100), .A2(n990), .ZN(n815) );
  NAND2_X1 U918 ( .A1(n816), .A2(n815), .ZN(n822) );
  NAND2_X1 U919 ( .A1(G112), .A2(n986), .ZN(n817) );
  XNOR2_X1 U920 ( .A(n817), .B(KEYINPUT106), .ZN(n820) );
  NAND2_X1 U921 ( .A1(G124), .A2(n985), .ZN(n818) );
  XNOR2_X1 U922 ( .A(n818), .B(KEYINPUT44), .ZN(n819) );
  NAND2_X1 U923 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U924 ( .A1(n822), .A2(n821), .ZN(G162) );
  XNOR2_X1 U925 ( .A(G16), .B(KEYINPUT56), .ZN(n848) );
  XNOR2_X1 U926 ( .A(G171), .B(G1961), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n949), .B(G1341), .ZN(n825) );
  XNOR2_X1 U928 ( .A(n823), .B(G1348), .ZN(n824) );
  NOR2_X1 U929 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U930 ( .A1(n827), .A2(n826), .ZN(n840) );
  XNOR2_X1 U931 ( .A(n828), .B(G1956), .ZN(n830) );
  NAND2_X1 U932 ( .A1(G1971), .A2(G303), .ZN(n829) );
  NAND2_X1 U933 ( .A1(n830), .A2(n829), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U935 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(KEYINPUT116), .B(n835), .Z(n836) );
  NOR2_X1 U937 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n838), .B(KEYINPUT117), .ZN(n839) );
  NOR2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(KEYINPUT118), .B(n841), .ZN(n846) );
  XNOR2_X1 U941 ( .A(G1966), .B(G168), .ZN(n843) );
  NAND2_X1 U942 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U943 ( .A(KEYINPUT57), .B(n844), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n880) );
  INV_X1 U946 ( .A(G16), .ZN(n878) );
  XNOR2_X1 U947 ( .A(G1986), .B(KEYINPUT124), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n849), .B(G24), .ZN(n855) );
  XNOR2_X1 U949 ( .A(G1976), .B(KEYINPUT122), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n850), .B(G23), .ZN(n852) );
  XNOR2_X1 U951 ( .A(G22), .B(G1971), .ZN(n851) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT123), .ZN(n854) );
  NOR2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U955 ( .A(KEYINPUT58), .B(n856), .ZN(n874) );
  XNOR2_X1 U956 ( .A(G1961), .B(G5), .ZN(n872) );
  XNOR2_X1 U957 ( .A(G1348), .B(KEYINPUT59), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(G4), .ZN(n862) );
  XOR2_X1 U959 ( .A(n858), .B(G20), .Z(n860) );
  XNOR2_X1 U960 ( .A(G6), .B(G1981), .ZN(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n865) );
  XOR2_X1 U963 ( .A(KEYINPUT119), .B(G1341), .Z(n863) );
  XNOR2_X1 U964 ( .A(G19), .B(n863), .ZN(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(n866), .B(KEYINPUT120), .Z(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT60), .B(n867), .ZN(n869) );
  XNOR2_X1 U968 ( .A(G21), .B(G1966), .ZN(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U970 ( .A(KEYINPUT121), .B(n870), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(KEYINPUT61), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT125), .B(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U976 ( .A1(n880), .A2(n879), .ZN(n904) );
  XOR2_X1 U977 ( .A(KEYINPUT55), .B(KEYINPUT114), .Z(n898) );
  XNOR2_X1 U978 ( .A(G2090), .B(G35), .ZN(n893) );
  XOR2_X1 U979 ( .A(G1991), .B(G25), .Z(n881) );
  NAND2_X1 U980 ( .A1(n881), .A2(G28), .ZN(n890) );
  XNOR2_X1 U981 ( .A(G1996), .B(G32), .ZN(n883) );
  XNOR2_X1 U982 ( .A(G33), .B(G2072), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n888) );
  XNOR2_X1 U984 ( .A(G2067), .B(G26), .ZN(n886) );
  XNOR2_X1 U985 ( .A(G27), .B(n884), .ZN(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(KEYINPUT53), .B(n891), .ZN(n892) );
  NOR2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n896) );
  XOR2_X1 U991 ( .A(G2084), .B(G34), .Z(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT54), .B(n894), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n900) );
  INV_X1 U995 ( .A(G29), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U997 ( .A1(G11), .A2(n901), .ZN(n902) );
  XOR2_X1 U998 ( .A(KEYINPUT115), .B(n902), .Z(n903) );
  NOR2_X1 U999 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n905), .B(KEYINPUT126), .ZN(n941) );
  INV_X1 U1001 ( .A(n906), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(n908), .A2(n907), .ZN(n933) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n989), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n990), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n917) );
  XNOR2_X1 U1006 ( .A(KEYINPUT108), .B(KEYINPUT47), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(n986), .A2(G115), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n985), .A2(G127), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT107), .B(n911), .Z(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n915), .B(n914), .Z(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n997) );
  XOR2_X1 U1013 ( .A(G2072), .B(n997), .Z(n919) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n921) );
  XOR2_X1 U1016 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n931) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n927) );
  NOR2_X1 U1023 ( .A1(n974), .A2(n927), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n936), .ZN(n938) );
  INV_X1 U1029 ( .A(KEYINPUT55), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(n939), .A2(G29), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1033 ( .A(KEYINPUT62), .B(n942), .Z(G311) );
  XNOR2_X1 U1034 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1035 ( .A(G120), .ZN(G236) );
  INV_X1 U1036 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(G325) );
  INV_X1 U1038 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1039 ( .A(KEYINPUT111), .B(n945), .Z(n948) );
  XNOR2_X1 U1040 ( .A(n946), .B(G286), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n948), .B(n947), .ZN(n951) );
  XOR2_X1 U1042 ( .A(n949), .B(G171), .Z(n950) );
  XNOR2_X1 U1043 ( .A(n951), .B(n950), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(G37), .A2(n952), .ZN(G397) );
  XOR2_X1 U1045 ( .A(G2096), .B(KEYINPUT43), .Z(n954) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G2072), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n954), .B(n953), .ZN(n955) );
  XOR2_X1 U1048 ( .A(n955), .B(KEYINPUT104), .Z(n957) );
  XNOR2_X1 U1049 ( .A(G2090), .B(G2678), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n957), .B(n956), .ZN(n961) );
  XOR2_X1 U1051 ( .A(KEYINPUT42), .B(G2100), .Z(n959) );
  XNOR2_X1 U1052 ( .A(G2078), .B(G2084), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n959), .B(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(G227) );
  XOR2_X1 U1055 ( .A(G2474), .B(G1971), .Z(n963) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G1966), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n963), .B(n962), .ZN(n967) );
  XOR2_X1 U1058 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n965) );
  XNOR2_X1 U1059 ( .A(G1991), .B(G1981), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n965), .B(n964), .ZN(n966) );
  XOR2_X1 U1061 ( .A(n967), .B(n966), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G1961), .B(G1976), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n971) );
  XOR2_X1 U1064 ( .A(G1986), .B(G1956), .Z(n970) );
  XNOR2_X1 U1065 ( .A(n971), .B(n970), .ZN(G229) );
  XOR2_X1 U1066 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(n973), .B(n972), .ZN(n978) );
  XOR2_X1 U1069 ( .A(G164), .B(n974), .Z(n975) );
  XNOR2_X1 U1070 ( .A(n976), .B(n975), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n978), .B(n977), .ZN(n984) );
  XOR2_X1 U1072 ( .A(G160), .B(G162), .Z(n979) );
  XNOR2_X1 U1073 ( .A(n980), .B(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n984), .B(n983), .ZN(n999) );
  NAND2_X1 U1076 ( .A1(G130), .A2(n985), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(G118), .A2(n986), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n995) );
  NAND2_X1 U1079 ( .A1(G142), .A2(n989), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(G106), .A2(n990), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1082 ( .A(KEYINPUT45), .B(n993), .Z(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n997), .B(n996), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n999), .B(n998), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(G37), .A2(n1000), .ZN(G395) );
  NOR2_X1 U1087 ( .A1(G227), .A2(G229), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT49), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(G397), .A2(n1002), .ZN(n1007) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(G401), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT112), .B(n1004), .Z(n1005) );
  NOR2_X1 U1092 ( .A1(G395), .A2(n1005), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(G225) );
  INV_X1 U1094 ( .A(G225), .ZN(G308) );
  INV_X1 U1095 ( .A(G108), .ZN(G238) );
endmodule

