//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  INV_X1    g002(.A(G131), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G137), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n194), .B1(new_n191), .B2(G137), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n192), .C1(new_n195), .C2(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n193), .A2(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n210), .A2(KEYINPUT64), .A3(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(new_n210), .B2(G146), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n207), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(G143), .B2(new_n206), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n210), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n206), .A2(G143), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n215), .A2(new_n208), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n196), .A2(new_n205), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n207), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n221), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n197), .A2(new_n199), .A3(G137), .ZN(new_n230));
  INV_X1    g044(.A(new_n194), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n190), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT11), .B1(new_n200), .B2(new_n201), .ZN(new_n233));
  OAI21_X1  g047(.A(G131), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n234), .B2(new_n196), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n188), .B1(new_n220), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n206), .B2(G143), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n210), .A2(KEYINPUT64), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n216), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n240), .A2(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(new_n231), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n189), .B1(new_n243), .B2(new_n192), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n232), .A2(new_n233), .A3(G131), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n219), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n213), .A2(new_n218), .A3(KEYINPUT67), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n196), .A3(new_n249), .A4(new_n205), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(KEYINPUT30), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G116), .ZN(new_n253));
  INV_X1    g067(.A(G116), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G119), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT2), .B(G113), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G113), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT2), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT2), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G113), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G116), .B(G119), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n265), .A3(KEYINPUT66), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n256), .A2(new_n257), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n236), .A2(new_n251), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n246), .A3(new_n250), .ZN(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT27), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n271), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n271), .A2(KEYINPUT31), .A3(new_n276), .A4(new_n281), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n270), .B1(new_n220), .B2(new_n235), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT28), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n276), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n281), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n284), .A2(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n187), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT72), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n289), .B1(new_n276), .B2(new_n286), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n213), .A2(KEYINPUT67), .A3(new_n218), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT67), .B1(new_n213), .B2(new_n218), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n189), .B1(new_n202), .B2(new_n203), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n232), .A2(new_n233), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(new_n189), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n234), .A2(new_n196), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n304), .A2(new_n307), .B1(new_n308), .B2(new_n241), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT28), .B1(new_n309), .B2(new_n275), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n301), .A2(new_n310), .A3(new_n292), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n311), .B2(KEYINPUT69), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n281), .B1(new_n271), .B2(new_n276), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n288), .A2(new_n281), .A3(new_n290), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  INV_X1    g134(.A(new_n274), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT68), .B1(new_n266), .B2(new_n268), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AND4_X1   g137(.A1(new_n248), .A2(new_n249), .A3(new_n196), .A4(new_n205), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n235), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n276), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n310), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n281), .A2(KEYINPUT29), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n320), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n289), .B1(new_n325), .B2(new_n276), .ZN(new_n331));
  NOR4_X1   g145(.A1(new_n331), .A2(new_n310), .A3(KEYINPUT71), .A4(new_n328), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n330), .A2(new_n332), .A3(G902), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n319), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G472), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n284), .A2(new_n285), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n291), .A2(new_n292), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n297), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n300), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT9), .B(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT77), .ZN(new_n343));
  INV_X1    g157(.A(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G221), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n346), .B(KEYINPUT78), .Z(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n215), .A2(new_n208), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n213), .B1(new_n240), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G104), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT3), .B1(new_n351), .B2(G107), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n353));
  INV_X1    g167(.A(G107), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(G104), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(G107), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n352), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n354), .A2(G104), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n351), .A2(G107), .ZN(new_n360));
  OAI21_X1  g174(.A(G101), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n348), .B1(new_n350), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n352), .A2(new_n355), .A3(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n367), .A3(G101), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(new_n369), .B2(new_n241), .ZN(new_n370));
  INV_X1    g184(.A(new_n308), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n358), .A2(new_n361), .A3(KEYINPUT10), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n304), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n248), .A2(new_n373), .A3(new_n372), .A4(new_n249), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n370), .B(new_n371), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n366), .A2(new_n241), .A3(new_n368), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n358), .A2(new_n361), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n228), .B1(new_n208), .B2(new_n215), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n213), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n380), .B1(new_n383), .B2(new_n348), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n248), .A2(new_n249), .A3(new_n373), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT80), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n386), .B2(new_n375), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT81), .A3(new_n371), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n379), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n387), .A2(new_n371), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G140), .ZN(new_n392));
  INV_X1    g206(.A(G953), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G227), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n392), .B(new_n394), .Z(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n350), .A2(new_n362), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n219), .B2(new_n362), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT12), .A3(new_n308), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n308), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT12), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n395), .B1(new_n379), .B2(new_n388), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g223(.A(KEYINPUT83), .B(new_n395), .C1(new_n379), .C2(new_n388), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n396), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n344), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n344), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n389), .A2(new_n406), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n415), .A2(new_n395), .B1(new_n407), .B2(new_n390), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n416), .B2(G469), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n347), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n252), .B2(G128), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n421), .B(new_n422), .C1(G119), .C2(new_n208), .ZN(new_n423));
  XNOR2_X1  g237(.A(G119), .B(G128), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT24), .B(G110), .Z(new_n425));
  AOI22_X1  g239(.A1(new_n423), .A2(G110), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G140), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G125), .ZN(new_n428));
  INV_X1    g242(.A(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G140), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT73), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(KEYINPUT73), .A3(G140), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT16), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT16), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n434), .A2(new_n206), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n206), .B1(new_n434), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n426), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G146), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n428), .A2(new_n430), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n206), .ZN(new_n443));
  OAI22_X1  g257(.A1(new_n423), .A2(G110), .B1(new_n424), .B2(new_n425), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n393), .A2(G221), .A3(G234), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT74), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G137), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n439), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n449), .B1(new_n439), .B2(new_n445), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT75), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n439), .A2(new_n445), .ZN(new_n454));
  INV_X1    g268(.A(new_n449), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT75), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(G234), .B2(new_n344), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G902), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n419), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  AOI211_X1 g278(.A(KEYINPUT76), .B(new_n464), .C1(new_n453), .C2(new_n458), .ZN(new_n465));
  INV_X1    g279(.A(new_n461), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n344), .A3(new_n450), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT25), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n456), .A2(KEYINPUT25), .A3(new_n344), .A4(new_n450), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n463), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n473));
  INV_X1    g287(.A(G237), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n393), .A3(G214), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n210), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n277), .A2(G143), .A3(G214), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT18), .A2(G131), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n432), .A2(G146), .A3(new_n433), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n443), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(G104), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT19), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n432), .B2(new_n433), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n442), .A2(KEYINPUT19), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n206), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n441), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n478), .B2(G131), .ZN(new_n494));
  AOI211_X1 g308(.A(KEYINPUT87), .B(new_n189), .C1(new_n476), .C2(new_n477), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n476), .A2(new_n189), .A3(new_n477), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n491), .A2(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n441), .A2(new_n490), .A3(KEYINPUT88), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n486), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n437), .A2(new_n438), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n475), .A2(new_n210), .ZN(new_n502));
  AOI21_X1  g316(.A(G143), .B1(new_n277), .B2(G214), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT87), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n478), .A2(new_n493), .A3(G131), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n497), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT17), .B1(new_n494), .B2(new_n495), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n501), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n485), .B1(new_n510), .B2(new_n483), .ZN(new_n511));
  NOR2_X1   g325(.A1(G475), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n500), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT20), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n473), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n483), .ZN(new_n517));
  INV_X1    g331(.A(new_n485), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n491), .A2(new_n492), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n496), .A2(new_n497), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n499), .ZN(new_n522));
  INV_X1    g336(.A(new_n486), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT89), .B(KEYINPUT20), .C1(new_n525), .C2(new_n513), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT20), .B1(new_n513), .B2(KEYINPUT90), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(KEYINPUT90), .B2(new_n513), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(KEYINPUT94), .A2(G952), .ZN(new_n531));
  NAND2_X1  g345(.A1(KEYINPUT94), .A2(G952), .ZN(new_n532));
  AOI21_X1  g346(.A(G953), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G234), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n474), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(G902), .B(G953), .C1(new_n534), .C2(new_n474), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT95), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT21), .B(G898), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n254), .A2(G122), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G122), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G116), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n545), .A3(new_n354), .ZN(new_n546));
  OAI21_X1  g360(.A(G107), .B1(new_n541), .B2(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n210), .A2(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n208), .A2(G143), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n191), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n210), .A2(KEYINPUT13), .A3(G128), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n553), .A2(new_n554), .A3(new_n550), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n548), .B(new_n551), .C1(new_n555), .C2(new_n193), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT14), .B1(new_n543), .B2(G116), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT92), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n541), .B1(new_n559), .B2(new_n544), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n354), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n551), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n191), .B1(new_n549), .B2(new_n550), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n546), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n556), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n343), .A2(G217), .A3(new_n393), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n556), .B(new_n566), .C1(new_n561), .C2(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n344), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n572), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n344), .A3(new_n569), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(KEYINPUT93), .A3(new_n575), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n540), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n517), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n344), .B1(new_n517), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g397(.A(G475), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n530), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G214), .B1(G237), .B2(G902), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n241), .A2(new_n429), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n219), .A2(G125), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n393), .A2(G224), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT85), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n366), .A2(new_n268), .A3(new_n266), .A4(new_n368), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT5), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n252), .A3(G116), .ZN(new_n595));
  OAI211_X1 g409(.A(G113), .B(new_n595), .C1(new_n256), .C2(new_n594), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n596), .A2(new_n265), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n362), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G122), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n593), .A2(new_n598), .A3(new_n600), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(KEYINPUT6), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT84), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT6), .ZN(new_n606));
  AND4_X1   g420(.A1(new_n605), .A2(new_n599), .A3(new_n606), .A4(new_n601), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n600), .B1(new_n593), .B2(new_n598), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n608), .B2(new_n606), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n592), .B(new_n604), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n597), .B1(KEYINPUT86), .B2(new_n381), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n596), .A2(new_n265), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT86), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n362), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n600), .B(KEYINPUT8), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n229), .A2(G125), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n617), .B(new_n619), .C1(G125), .C2(new_n219), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n618), .B1(new_n587), .B2(new_n588), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n622), .B2(new_n603), .ZN(new_n623));
  OAI21_X1  g437(.A(G210), .B1(G237), .B2(G902), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n610), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n610), .B2(new_n623), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n586), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n585), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n341), .A2(new_n418), .A3(new_n472), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  OAI21_X1  g444(.A(G472), .B1(new_n293), .B2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n338), .A2(new_n294), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n418), .A2(new_n472), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(KEYINPUT96), .B(new_n586), .C1(new_n625), .C2(new_n626), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n540), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n566), .A2(KEYINPUT98), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n565), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n565), .B2(new_n641), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n568), .A2(new_n569), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n571), .A2(G902), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n646), .A2(new_n647), .B1(new_n571), .B2(new_n570), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n530), .B2(new_n584), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n638), .A2(new_n639), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n634), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND2_X1  g467(.A1(new_n514), .A2(new_n515), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n516), .A2(new_n526), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n578), .A2(new_n579), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n584), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n540), .B(new_n657), .C1(new_n636), .C2(new_n637), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n634), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT99), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT100), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n413), .A2(new_n417), .ZN(new_n665));
  INV_X1    g479(.A(new_n347), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n455), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n454), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n464), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n471), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n585), .A2(new_n627), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n665), .A2(new_n666), .A3(new_n672), .A4(new_n633), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AND3_X1   g489(.A1(new_n340), .A2(new_n296), .A3(new_n299), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n671), .B1(new_n676), .B2(new_n335), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n536), .B1(new_n678), .B2(new_n538), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n638), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n677), .A2(new_n418), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n530), .A2(new_n584), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n684), .A2(new_n656), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n586), .A3(new_n671), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n610), .A2(new_n623), .ZN(new_n690));
  INV_X1    g504(.A(new_n624), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n610), .A2(new_n623), .A3(new_n624), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n326), .A2(new_n292), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n282), .A2(new_n697), .A3(KEYINPUT101), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n344), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT101), .B1(new_n282), .B2(new_n697), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n676), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n679), .B(KEYINPUT39), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n418), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n696), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(KEYINPUT40), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  AOI211_X1 g523(.A(new_n648), .B(new_n679), .C1(new_n530), .C2(new_n584), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n638), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT104), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n638), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n677), .A2(new_n712), .A3(new_n418), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  INV_X1    g530(.A(new_n472), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n676), .B2(new_n335), .ZN(new_n718));
  INV_X1    g532(.A(new_n650), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n411), .A2(new_n412), .A3(new_n344), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n412), .B1(new_n411), .B2(new_n344), .ZN(new_n721));
  INV_X1    g535(.A(new_n346), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n719), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND3_X1  g540(.A1(new_n718), .A2(new_n723), .A3(new_n658), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT105), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n723), .A3(new_n729), .A4(new_n658), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  INV_X1    g546(.A(new_n585), .ZN(new_n733));
  INV_X1    g547(.A(new_n671), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n340), .A2(new_n296), .A3(new_n299), .ZN(new_n735));
  INV_X1    g549(.A(G472), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n319), .B2(new_n333), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n395), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n389), .B2(new_n390), .ZN(new_n740));
  INV_X1    g554(.A(new_n406), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n377), .A2(new_n378), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT81), .B1(new_n387), .B2(new_n371), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n744), .B2(KEYINPUT83), .ZN(new_n745));
  INV_X1    g559(.A(new_n410), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(G469), .B1(new_n747), .B2(G902), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n638), .A3(new_n346), .A4(new_n413), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n252), .ZN(G21));
  OAI21_X1  g565(.A(new_n292), .B1(new_n331), .B2(new_n310), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n336), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n294), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n631), .A2(new_n754), .A3(new_n472), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n639), .A3(new_n638), .A4(new_n685), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n748), .A2(new_n346), .A3(new_n413), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n543), .ZN(G24));
  INV_X1    g573(.A(new_n749), .ZN(new_n760));
  INV_X1    g574(.A(new_n679), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n649), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n631), .A2(new_n754), .A3(new_n734), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NOR2_X1   g580(.A1(new_n625), .A2(new_n626), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n586), .A3(new_n346), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n413), .B2(new_n417), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n341), .A2(new_n769), .A3(new_n472), .A4(new_n710), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n338), .A2(new_n297), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n296), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT106), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n296), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n335), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n762), .A2(new_n771), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n472), .A3(new_n769), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n772), .A2(KEYINPUT107), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n189), .ZN(G33));
  NAND4_X1  g600(.A1(new_n341), .A2(new_n769), .A3(new_n472), .A4(new_n680), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  INV_X1    g602(.A(new_n648), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n530), .A3(new_n584), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT43), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n633), .A2(new_n671), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(KEYINPUT44), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n767), .A2(new_n586), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  INV_X1    g618(.A(new_n416), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n412), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n416), .A2(KEYINPUT45), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n414), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT46), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n720), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n414), .B1(new_n807), .B2(new_n808), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n722), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n704), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n803), .A2(new_n804), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(KEYINPUT47), .ZN(new_n821));
  INV_X1    g635(.A(new_n815), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n413), .B1(new_n814), .B2(KEYINPUT46), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n346), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n800), .A2(new_n717), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n341), .A2(new_n828), .A3(new_n762), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n820), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n829), .ZN(new_n831));
  AOI211_X1 g645(.A(KEYINPUT110), .B(new_n831), .C1(new_n821), .C2(new_n826), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  NAND2_X1  g648(.A1(new_n793), .A2(new_n536), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT115), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n757), .A2(new_n799), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT48), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n472), .A3(new_n778), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(KEYINPUT48), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n841), .B(new_n842), .Z(new_n843));
  AND2_X1   g657(.A1(new_n836), .A2(new_n755), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n760), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n703), .A2(new_n472), .A3(new_n536), .A4(new_n837), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n684), .A2(new_n789), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n845), .A2(new_n533), .A3(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n846), .A2(new_n684), .A3(new_n789), .ZN(new_n850));
  INV_X1    g664(.A(new_n763), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n757), .A2(new_n586), .A3(new_n695), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT116), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n844), .A2(KEYINPUT50), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT50), .B1(new_n844), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n720), .A2(new_n721), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n666), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n844), .B(new_n800), .C1(new_n827), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n843), .B(new_n849), .C1(new_n857), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n857), .A2(new_n864), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n472), .B1(new_n735), .B2(new_n737), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n757), .A2(new_n870), .A3(new_n650), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n750), .A3(new_n758), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n694), .A2(new_n586), .A3(new_n639), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n530), .A2(new_n576), .A3(new_n584), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n847), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n876), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n634), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n418), .A2(new_n628), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n673), .B1(new_n881), .B2(new_n870), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n655), .A2(new_n584), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n799), .A2(new_n884), .A3(new_n576), .A4(new_n679), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n341), .A2(new_n418), .A3(new_n734), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n764), .A2(new_n769), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n886), .A2(new_n787), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n731), .A2(new_n872), .A3(new_n883), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT112), .B1(new_n785), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n772), .A2(KEYINPUT107), .A3(new_n780), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT107), .B1(new_n772), .B2(new_n780), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n738), .A2(new_n749), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n638), .A2(new_n685), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n723), .A2(new_n639), .A3(new_n896), .A4(new_n755), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n897), .A3(new_n724), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n730), .B2(new_n728), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n629), .B(new_n673), .C1(new_n634), .C2(new_n879), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n787), .A3(new_n887), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n893), .A2(new_n894), .A3(new_n899), .A4(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n890), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n734), .B2(new_n679), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n671), .A2(KEYINPUT113), .A3(new_n761), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n722), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n896), .A2(new_n702), .A3(new_n665), .A4(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n715), .A2(new_n765), .A3(new_n682), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT52), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n418), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n638), .A2(new_n713), .A3(new_n710), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n713), .B1(new_n638), .B2(new_n710), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n919), .B2(new_n681), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(KEYINPUT52), .A3(new_n765), .A4(new_n910), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n913), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n913), .A2(new_n922), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n913), .A2(new_n921), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n890), .A2(new_n903), .A3(new_n926), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n905), .A2(new_n925), .B1(KEYINPUT53), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n904), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n904), .B1(new_n772), .B2(new_n780), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n902), .A2(new_n731), .A3(new_n872), .A4(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n923), .A2(new_n924), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(KEYINPUT54), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n869), .A2(new_n929), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(G952), .B2(G953), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n472), .A2(new_n586), .A3(new_n666), .ZN(new_n939));
  OR3_X1    g753(.A1(new_n695), .A2(new_n790), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(KEYINPUT49), .B2(new_n859), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n703), .C1(KEYINPUT49), .C2(new_n859), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n938), .A2(new_n942), .ZN(G75));
  NOR2_X1   g757(.A1(new_n393), .A2(G952), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n935), .A2(new_n945), .A3(G902), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n933), .B1(new_n927), .B2(new_n904), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT120), .B1(new_n947), .B2(new_n344), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n691), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(new_n592), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(KEYINPUT56), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n944), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT119), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n935), .A2(G210), .A3(G902), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n955), .B1(new_n958), .B2(new_n952), .ZN(new_n959));
  INV_X1    g773(.A(new_n952), .ZN(new_n960));
  AOI211_X1 g774(.A(KEYINPUT119), .B(new_n960), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n954), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT121), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT121), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n954), .B(new_n964), .C1(new_n959), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(G51));
  XNOR2_X1  g780(.A(new_n935), .B(KEYINPUT54), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n414), .B(KEYINPUT57), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n411), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n946), .A2(new_n948), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(new_n809), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n944), .B1(new_n970), .B2(new_n972), .ZN(G54));
  NAND2_X1  g787(.A1(KEYINPUT58), .A2(G475), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n525), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n944), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n971), .A2(new_n525), .A3(new_n974), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(G60));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n936), .B2(new_n929), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT122), .B1(new_n982), .B2(new_n646), .ZN(new_n983));
  INV_X1    g797(.A(new_n646), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n981), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n944), .B1(new_n967), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n982), .A2(KEYINPUT122), .A3(new_n646), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G63));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT60), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n935), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n453), .A3(new_n458), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n976), .C1(new_n669), .C2(new_n992), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT61), .Z(G66));
  INV_X1    g809(.A(G224), .ZN(new_n996));
  OAI21_X1  g810(.A(G953), .B1(new_n539), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n899), .A2(new_n883), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n997), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n950), .B1(G898), .B2(new_n393), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  AND2_X1   g816(.A1(new_n920), .A2(new_n765), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n708), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT62), .Z(new_n1005));
  OAI21_X1  g819(.A(new_n818), .B1(new_n830), .B2(new_n832), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n718), .B(new_n800), .C1(new_n877), .C2(new_n878), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n1005), .B(new_n1007), .C1(new_n705), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n393), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n236), .A2(new_n251), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n488), .A2(new_n489), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  XOR2_X1   g827(.A(KEYINPUT123), .B(KEYINPUT124), .Z(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n817), .A2(new_n472), .A3(new_n896), .A4(new_n778), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1017), .A2(new_n893), .A3(new_n787), .A4(new_n1003), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1019), .A2(new_n833), .A3(KEYINPUT125), .A4(new_n818), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT125), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1021), .B1(new_n1006), .B2(new_n1018), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n1022), .A3(new_n393), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1015), .B1(G900), .B2(G953), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n393), .B1(G227), .B2(G900), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1026), .B(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n1009), .B2(new_n998), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n271), .A2(new_n276), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1031), .A2(new_n1032), .A3(new_n281), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n314), .A2(new_n315), .A3(new_n282), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n928), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1020), .A2(new_n1022), .A3(new_n999), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1037), .A2(new_n1038), .A3(new_n1030), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1032), .A2(new_n281), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1038), .B1(new_n1037), .B2(new_n1030), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n976), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT127), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT127), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1045), .B(new_n976), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1036), .B1(new_n1044), .B2(new_n1046), .ZN(G57));
endmodule


