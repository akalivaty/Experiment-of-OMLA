//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G101), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(KEYINPUT68), .B(KEYINPUT3), .C1(new_n461), .C2(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT67), .Z(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(G2104), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n462), .A2(new_n465), .A3(new_n468), .A4(new_n472), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n472), .B2(G112), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n462), .A2(new_n465), .A3(new_n468), .A4(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G124), .ZN(G162));
  NAND4_X1  g064(.A1(new_n476), .A2(new_n477), .A3(G138), .A4(new_n472), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n482), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n487), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n494), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT5), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n501), .A2(new_n504), .B1(new_n500), .B2(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(new_n503), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(new_n511), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(G63), .A2(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n512), .A2(G51), .B1(new_n505), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n520), .B(new_n523), .C1(new_n524), .C2(new_n515), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(G651), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n501), .A2(new_n504), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n500), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n511), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT74), .B(G52), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n537), .A2(G90), .B1(new_n512), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n507), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n512), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n515), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n512), .A2(new_n554), .A3(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n534), .A2(G65), .A3(new_n535), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT76), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n561), .B(new_n558), .C1(new_n536), .C2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n563), .A3(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n537), .A2(G91), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  OAI21_X1  g143(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n537), .A2(G87), .B1(G49), .B2(new_n512), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AND3_X1   g148(.A1(new_n505), .A2(G86), .A3(new_n514), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT79), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n512), .A2(G48), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n536), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n505), .A2(KEYINPUT78), .A3(G61), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n575), .A2(new_n576), .A3(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n507), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n512), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n515), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  AOI22_X1  g166(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n507), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n596), .A2(G54), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT10), .B1(new_n515), .B2(new_n594), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n593), .A2(new_n595), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n601), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G168), .B2(new_n601), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(G168), .B2(new_n601), .ZN(G280));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  INV_X1    g185(.A(new_n547), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n601), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n600), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n601), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n617), .B(new_n618), .C1(G111), .C2(new_n472), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n482), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n488), .B2(G123), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n467), .A2(new_n461), .A3(G2105), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT13), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT83), .Z(G156));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  OAI21_X1  g208(.A(KEYINPUT14), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT85), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n638), .B(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(G14), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT86), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n651), .B(KEYINPUT17), .Z(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(new_n649), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n649), .A3(new_n647), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n650), .A2(new_n651), .A3(new_n647), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n664), .A3(new_n667), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n673), .C1(new_n664), .C2(new_n672), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n674), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT88), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  INV_X1    g258(.A(G288), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT33), .ZN(new_n686));
  INV_X1    g261(.A(G1976), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(G166), .A2(new_n682), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n682), .B2(G22), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n688), .A2(new_n689), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n682), .A2(G6), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G305), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT32), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n696), .A2(KEYINPUT34), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n695), .B2(new_n701), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G25), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n488), .A2(G119), .ZN(new_n709));
  INV_X1    g284(.A(G131), .ZN(new_n710));
  NOR2_X1   g285(.A1(G95), .A2(G2105), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n482), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT89), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n715), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n682), .A2(G24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n590), .B2(new_n682), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1986), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n706), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G141), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n482), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G129), .B2(new_n488), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n461), .A2(G2105), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G105), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G32), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  NOR2_X1   g315(.A1(G164), .A2(new_n707), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G27), .B2(new_n707), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n707), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT95), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  INV_X1    g321(.A(G140), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n482), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(G104), .A2(G2105), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n748), .B(new_n751), .C1(G128), .C2(new_n488), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(new_n707), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n753), .A2(new_n754), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n746), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  AND2_X1   g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  NOR2_X1   g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n707), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n763), .B(new_n764), .C1(new_n480), .C2(new_n707), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT99), .ZN(new_n769));
  OR4_X1    g344(.A1(new_n743), .A2(new_n759), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G21), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G168), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G35), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G162), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT29), .B(G2090), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n608), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n682), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n547), .B2(new_n682), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT92), .B(G1341), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G28), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n792), .A2(new_n793), .A3(new_n707), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n622), .A2(G29), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n786), .A2(new_n790), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n770), .A2(new_n779), .A3(new_n785), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n706), .B(new_n725), .C1(KEYINPUT91), .C2(KEYINPUT36), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n682), .A2(G5), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G171), .B2(new_n682), .ZN(new_n800));
  INV_X1    g375(.A(G1961), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n728), .A2(new_n797), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n476), .A2(new_n477), .A3(G127), .ZN(new_n804));
  INV_X1    g379(.A(G115), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n461), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G2105), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT96), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n732), .A2(G103), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT25), .Z(new_n810));
  INV_X1    g385(.A(G139), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n810), .C1(new_n811), .C2(new_n482), .ZN(new_n812));
  MUX2_X1   g387(.A(G33), .B(new_n812), .S(G29), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2072), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n682), .A2(KEYINPUT23), .A3(G20), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n816));
  INV_X1    g391(.A(G20), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n815), .B(new_n818), .C1(new_n819), .C2(new_n682), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT100), .B(G1956), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT101), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n803), .A2(new_n814), .A3(new_n824), .ZN(G311));
  OR3_X1    g400(.A1(new_n803), .A2(new_n814), .A3(new_n824), .ZN(G150));
  NAND2_X1  g401(.A1(new_n608), .A2(G559), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT39), .Z(new_n828));
  AOI22_X1  g403(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n507), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n512), .A2(G55), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n515), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n547), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n828), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT102), .B(G860), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT103), .Z(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n830), .B2(new_n833), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  INV_X1    g418(.A(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n482), .A2(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n488), .B2(G130), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n714), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n498), .A2(KEYINPUT104), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n851), .B(new_n496), .C1(new_n487), .C2(new_n497), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n494), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n849), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n812), .B(new_n626), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n752), .B(KEYINPUT105), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n737), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n622), .B(G160), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(G162), .Z(new_n863));
  OR3_X1    g438(.A1(new_n861), .A2(KEYINPUT106), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT106), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g443(.A1(new_n819), .A2(new_n600), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n608), .A2(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT107), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n869), .A2(new_n870), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n874), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n877), .B2(new_n872), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n835), .B(new_n613), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT108), .B1(new_n879), .B2(new_n876), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n880), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n886), .B(new_n887), .C1(new_n881), .C2(new_n882), .ZN(new_n888));
  XNOR2_X1  g463(.A(G166), .B(KEYINPUT109), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(G290), .B(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n885), .B2(new_n888), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n834), .A2(G868), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G295));
  NAND2_X1  g474(.A1(new_n885), .A2(new_n888), .ZN(new_n900));
  INV_X1    g475(.A(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n601), .B1(new_n902), .B2(new_n893), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT110), .B1(new_n903), .B2(new_n897), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n896), .A2(new_n905), .A3(new_n898), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(G331));
  XNOR2_X1  g482(.A(G168), .B(G171), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n835), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(KEYINPUT41), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n877), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(new_n892), .C1(new_n871), .C2(new_n910), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n878), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n871), .B2(new_n909), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n914), .B2(new_n901), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n914), .A2(new_n901), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT43), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n917), .A3(new_n915), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n919), .A2(new_n915), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n917), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n925), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g501(.A(KEYINPUT126), .ZN(new_n927));
  OR2_X1    g502(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n928));
  NAND2_X1  g503(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n819), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n855), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n473), .A2(G40), .A3(new_n479), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n494), .B2(new_n498), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT56), .B(G2072), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n494), .B1(new_n850), .B2(new_n852), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT50), .B1(new_n942), .B2(G1384), .ZN(new_n943));
  INV_X1    g518(.A(new_n937), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G1956), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n932), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1956), .ZN(new_n949));
  INV_X1    g524(.A(new_n943), .ZN(new_n950));
  INV_X1    g525(.A(new_n935), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(KEYINPUT50), .B2(new_n937), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(new_n930), .A3(new_n931), .A4(new_n940), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n942), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n782), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT119), .ZN(new_n959));
  NOR4_X1   g534(.A1(new_n942), .A2(new_n935), .A3(G1384), .A4(G2067), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n855), .A2(new_n945), .A3(new_n933), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n935), .B1(KEYINPUT50), .B2(new_n937), .ZN(new_n964));
  AOI21_X1  g539(.A(G1348), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT119), .B1(new_n965), .B2(new_n960), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n954), .A2(new_n608), .A3(new_n962), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1996), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n934), .A2(new_n968), .A3(new_n938), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT120), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n853), .B2(new_n854), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n951), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT58), .B(G1341), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n934), .A2(KEYINPUT120), .A3(new_n968), .A4(new_n938), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n547), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n977), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n547), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT122), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n948), .A2(new_n954), .A3(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n948), .B2(new_n954), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n980), .B(new_n981), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n965), .A2(KEYINPUT119), .A3(new_n960), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n959), .B1(new_n958), .B2(new_n961), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT60), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT60), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n966), .A2(new_n962), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n608), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT60), .B(new_n600), .C1(new_n988), .C2(new_n989), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n948), .B(new_n967), .C1(new_n987), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n855), .A2(new_n933), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n935), .B1(new_n997), .B2(new_n936), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT125), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n740), .A2(KEYINPUT53), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n934), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n936), .B1(new_n942), .B2(G1384), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n934), .A2(new_n1002), .A3(new_n951), .A4(new_n1000), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n934), .A2(new_n740), .A3(new_n938), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1007));
  NAND2_X1  g582(.A1(new_n963), .A2(new_n964), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1006), .A2(new_n1007), .B1(new_n1008), .B2(new_n801), .ZN(new_n1009));
  AOI21_X1  g584(.A(G301), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n944), .A2(KEYINPUT45), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n998), .A2(new_n1011), .A3(new_n1000), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n801), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G171), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1010), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT115), .B(G8), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1002), .A2(new_n951), .A3(new_n1011), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n773), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n963), .A2(new_n766), .A3(new_n964), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1019), .B(new_n1020), .C1(new_n1024), .C2(G286), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1020), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G168), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n1019), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n955), .A2(new_n957), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n766), .A2(new_n1029), .B1(new_n1021), .B2(new_n773), .ZN(new_n1030));
  INV_X1    g605(.A(G8), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1025), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1035));
  NAND3_X1  g610(.A1(new_n1005), .A2(G301), .A3(new_n1009), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1015), .A2(G171), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1018), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n942), .A2(new_n936), .A3(G1384), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n937), .A2(new_n936), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n951), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n692), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT111), .B(new_n692), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n963), .A2(new_n1048), .A3(new_n964), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT112), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n963), .A2(new_n1051), .A3(new_n1048), .A4(new_n964), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(new_n1053), .A3(KEYINPUT113), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1056), .A2(G8), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n574), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n583), .A2(new_n576), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G1981), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT116), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n575), .A2(new_n700), .A3(new_n583), .A4(new_n576), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(new_n1068), .A3(G1981), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n973), .A2(new_n1020), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1066), .A2(KEYINPUT49), .A3(new_n1069), .A4(new_n1067), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(G1976), .B2(new_n684), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1077), .B(new_n1078), .C1(G1976), .C2(new_n684), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n950), .A2(G2090), .A3(new_n952), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1043), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1020), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1059), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1062), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n996), .A2(new_n1039), .A3(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1030), .A2(G286), .A3(new_n1026), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1062), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1081), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1076), .A2(new_n687), .A3(new_n684), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1067), .B(KEYINPUT117), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1074), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1076), .A2(new_n1079), .A3(new_n1088), .A4(new_n1080), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1056), .A2(G8), .A3(new_n1061), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1059), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1092), .B(new_n1096), .C1(new_n1089), .C2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n927), .B1(new_n1087), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1037), .B1(new_n1034), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1086), .B(new_n1103), .C1(new_n1102), .C2(new_n1034), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1059), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n1081), .A3(new_n1088), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1106), .A2(KEYINPUT63), .B1(new_n1074), .B2(new_n1095), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n996), .A2(new_n1086), .A3(new_n1039), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(KEYINPUT126), .A4(new_n1092), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1101), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1002), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n951), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G2067), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n752), .B(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n737), .B(G1996), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n717), .B1(new_n709), .B2(new_n713), .ZN(new_n1118));
  OR3_X1    g693(.A1(new_n709), .A2(new_n713), .A3(new_n717), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1986), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n590), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G290), .A2(G1986), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1113), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1110), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1113), .B1(new_n1115), .B2(new_n737), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1113), .A2(KEYINPUT46), .A3(new_n968), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT46), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1112), .B2(G1996), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT127), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT47), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n752), .A2(new_n1114), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1117), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1113), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1113), .A2(new_n1123), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT48), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1132), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1125), .A2(new_n1140), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g716(.A1(G401), .A2(G229), .ZN(new_n1143));
  INV_X1    g717(.A(new_n922), .ZN(new_n1144));
  AOI21_X1  g718(.A(new_n917), .B1(new_n919), .B2(new_n915), .ZN(new_n1145));
  OAI211_X1 g719(.A(new_n661), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g720(.A1(new_n867), .A2(G319), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1147), .ZN(G308));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1149));
  NAND4_X1  g723(.A1(new_n1149), .A2(new_n924), .A3(new_n661), .A4(new_n1143), .ZN(G225));
endmodule


