//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  OR2_X1    g000(.A1(KEYINPUT66), .A2(G116), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT66), .A2(G116), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G119), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT2), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n192), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n189), .B2(new_n192), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n203), .A2(KEYINPUT3), .A3(G107), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(KEYINPUT80), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G104), .ZN(new_n208));
  AOI21_X1  g022(.A(G107), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n205), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT80), .B(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(G101), .B(new_n202), .C1(new_n211), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n208), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n204), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n220), .B2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n216), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT4), .B1(new_n211), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n201), .B(new_n215), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n225), .A2(new_n216), .A3(new_n205), .A4(new_n213), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n218), .A2(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n209), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n189), .A2(KEYINPUT5), .A3(new_n192), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n193), .B1(new_n191), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n228), .A3(new_n232), .A4(new_n198), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n233), .A3(new_n235), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G953), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT64), .B(G128), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(G143), .B2(new_n241), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n242), .A2(new_n244), .A3(new_n247), .A4(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(G125), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  OR2_X1    g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n245), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n242), .A2(new_n244), .A3(new_n254), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(G224), .B(new_n240), .C1(new_n251), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n240), .A2(G224), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n242), .A2(new_n244), .B1(new_n253), .B2(new_n254), .ZN(new_n261));
  INV_X1    g075(.A(new_n257), .ZN(new_n262));
  OAI21_X1  g076(.A(G125), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT64), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n268), .A2(new_n269), .B1(new_n242), .B2(new_n244), .ZN(new_n270));
  INV_X1    g084(.A(new_n250), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n260), .B(new_n263), .C1(new_n272), .C2(G125), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n259), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n234), .A2(new_n275), .A3(new_n236), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n239), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n235), .B(KEYINPUT8), .ZN(new_n280));
  AND4_X1   g094(.A1(new_n226), .A2(new_n228), .A3(new_n198), .A4(new_n232), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n226), .A2(new_n228), .B1(new_n232), .B2(new_n198), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT7), .B1(new_n240), .B2(G224), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n259), .B2(new_n273), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(new_n260), .C1(new_n251), .C2(new_n258), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n283), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n224), .A2(new_n233), .A3(new_n235), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n278), .B(new_n279), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n238), .B(new_n283), .C1(new_n285), .C2(new_n288), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n278), .B1(new_n293), .B2(new_n279), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n296), .B(new_n277), .C1(new_n292), .C2(new_n294), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n279), .B1(new_n289), .B2(new_n290), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT85), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n291), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n304), .B2(new_n277), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT86), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  INV_X1    g122(.A(G217), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n308), .A2(new_n309), .A3(G953), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT14), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n187), .A2(G122), .A3(new_n188), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT89), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT89), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n187), .A2(new_n314), .A3(G122), .A4(new_n188), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n190), .A2(G122), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT91), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT66), .A2(G116), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT66), .A2(G116), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n321), .B2(G122), .ZN(new_n322));
  INV_X1    g136(.A(G122), .ZN(new_n323));
  NOR4_X1   g137(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT89), .A4(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT14), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n326));
  INV_X1    g140(.A(new_n317), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n313), .A2(new_n311), .A3(new_n315), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n318), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G107), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n246), .A2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n243), .A2(G128), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G134), .ZN(new_n335));
  INV_X1    g149(.A(G134), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n336), .A3(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n313), .A2(new_n315), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n218), .A3(new_n327), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n327), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G107), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n340), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT13), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n246), .A2(G143), .B1(new_n347), .B2(new_n333), .ZN(new_n348));
  INV_X1    g162(.A(new_n333), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT90), .B1(new_n349), .B2(KEYINPUT13), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n352));
  OAI21_X1  g166(.A(G134), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n346), .B(new_n337), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n310), .B1(new_n343), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n341), .B1(new_n330), .B2(G107), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n337), .B1(new_n351), .B2(new_n353), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n340), .B2(new_n345), .ZN(new_n358));
  INV_X1    g172(.A(new_n310), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n279), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G478), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT94), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n329), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n325), .A2(new_n327), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(KEYINPUT91), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n218), .B1(new_n370), .B2(new_n328), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n354), .B(new_n310), .C1(new_n371), .C2(new_n341), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n359), .B1(new_n356), .B2(new_n358), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n375));
  INV_X1    g189(.A(new_n366), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n361), .A2(KEYINPUT93), .A3(new_n366), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n374), .B2(new_n376), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT16), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n252), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n384), .A2(G146), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G146), .B1(new_n384), .B2(new_n385), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n240), .A3(G214), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n243), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT17), .A3(G131), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT87), .B1(new_n391), .B2(G131), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(G131), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n390), .B(G143), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n396));
  INV_X1    g210(.A(G131), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n388), .B(new_n392), .C1(new_n399), .C2(KEYINPUT17), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n203), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n395), .B1(new_n403), .B2(new_n397), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n383), .B(new_n241), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n383), .B(KEYINPUT19), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n386), .B1(new_n241), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n399), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n407), .ZN(new_n412));
  INV_X1    g226(.A(new_n402), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(G475), .A2(G902), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT88), .B1(new_n408), .B2(new_n414), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(KEYINPUT20), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(KEYINPUT88), .A3(new_n420), .A4(new_n416), .ZN(new_n421));
  INV_X1    g235(.A(new_n408), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n402), .B1(new_n400), .B2(new_n407), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n279), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n419), .A2(new_n421), .B1(G475), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n378), .A2(new_n382), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G952), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n428), .A2(KEYINPUT95), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(KEYINPUT95), .ZN(new_n430));
  AOI21_X1  g244(.A(G953), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G234), .A2(G237), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n432), .A2(G902), .A3(G953), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G214), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n307), .A2(new_n427), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n240), .A2(G227), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT79), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G140), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n336), .B2(G137), .ZN(new_n449));
  INV_X1    g263(.A(G137), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT11), .A3(G134), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n336), .A2(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n451), .A3(new_n397), .A4(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n245), .B1(new_n248), .B2(new_n264), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n250), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n226), .A2(new_n228), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n249), .A2(new_n250), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n226), .B2(new_n228), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI211_X1 g277(.A(KEYINPUT83), .B(new_n460), .C1(new_n226), .C2(new_n228), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n456), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT12), .B(new_n456), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n226), .A2(new_n228), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n272), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n470), .A2(new_n472), .B1(new_n459), .B2(new_n471), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n256), .A2(new_n257), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n215), .C1(new_n221), .C2(new_n223), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n456), .B(KEYINPUT82), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n469), .A2(KEYINPUT84), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT84), .B1(new_n469), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n447), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n477), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(new_n447), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(new_n475), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n456), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(G469), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G469), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n279), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n482), .A2(new_n469), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n477), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n447), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n443), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT69), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n389), .A2(new_n240), .A3(G210), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT68), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(KEYINPUT68), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n500), .A2(new_n505), .B1(new_n503), .B2(new_n502), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n496), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT69), .A3(new_n506), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n199), .A2(new_n200), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n336), .A2(G137), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n450), .A2(G134), .ZN(new_n516));
  OAI21_X1  g330(.A(G131), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n455), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n474), .A2(new_n456), .B1(new_n518), .B2(new_n460), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n456), .A2(new_n474), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n460), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT70), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n513), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n522), .A2(new_n514), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT28), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n512), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n514), .B1(new_n519), .B2(KEYINPUT30), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT65), .B(KEYINPUT30), .C1(new_n522), .C2(new_n523), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n514), .A3(new_n523), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n510), .A2(new_n506), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT31), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT65), .B1(new_n519), .B2(KEYINPUT30), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n524), .A2(new_n532), .A3(new_n533), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n527), .B1(new_n545), .B2(new_n531), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n539), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n530), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n495), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n530), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT31), .B1(new_n546), .B2(new_n539), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n201), .B1(new_n524), .B2(new_n533), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n544), .B2(new_n543), .ZN(new_n555));
  NOR4_X1   g369(.A1(new_n555), .A2(new_n541), .A3(new_n527), .A4(new_n538), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n552), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT32), .A3(new_n549), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n526), .A2(KEYINPUT72), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n455), .A2(new_n517), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n249), .B2(new_n250), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n454), .A2(new_n455), .B1(new_n256), .B2(new_n257), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n201), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n564), .B2(new_n537), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT28), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n568), .B(new_n513), .C1(new_n521), .C2(new_n525), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n538), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n559), .A2(new_n567), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n539), .B1(new_n536), .B2(new_n537), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n529), .A2(new_n512), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n201), .B1(new_n524), .B2(KEYINPUT70), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n519), .A2(new_n520), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT28), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n570), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n572), .B(new_n279), .C1(new_n573), .C2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n579), .A2(new_n580), .A3(G472), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n579), .B2(G472), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n551), .B(new_n558), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n309), .B1(G234), .B2(new_n279), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT78), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n240), .A2(G221), .A3(G234), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT77), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n587), .B(new_n589), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G119), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G128), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n268), .B2(new_n596), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT24), .B(G110), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT75), .B1(new_n596), .B2(G128), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n596), .A2(KEYINPUT75), .A3(G128), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT23), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(KEYINPUT74), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(KEYINPUT74), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n601), .B(new_n602), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n246), .A2(KEYINPUT23), .A3(G119), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n600), .B1(new_n608), .B2(G110), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n383), .A2(new_n241), .ZN(new_n610));
  INV_X1    g424(.A(new_n386), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI22_X1  g427(.A1(new_n386), .A2(new_n387), .B1(new_n598), .B2(new_n599), .ZN(new_n614));
  INV_X1    g428(.A(G110), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT76), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n608), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n606), .A2(KEYINPUT76), .A3(new_n607), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n595), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n612), .B(new_n593), .C1(new_n621), .C2(new_n614), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n622), .A3(new_n279), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n584), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n620), .A2(new_n622), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n584), .A2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n494), .A2(new_n583), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n441), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n216), .ZN(G3));
  INV_X1    g449(.A(new_n437), .ZN(new_n636));
  INV_X1    g450(.A(new_n300), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n438), .B(new_n636), .C1(new_n637), .C2(new_n305), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n362), .A2(G902), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT33), .B1(new_n355), .B2(new_n360), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n372), .A2(new_n373), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n374), .A2(G478), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n372), .A2(new_n373), .A3(new_n645), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n645), .B1(new_n372), .B2(new_n373), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n642), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n361), .A2(new_n362), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(KEYINPUT97), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n425), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n640), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI211_X1 g471(.A(KEYINPUT98), .B(new_n425), .C1(new_n649), .C2(new_n654), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n639), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n557), .B2(new_n279), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT96), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n548), .A2(new_n550), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n548), .B2(G902), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT96), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n494), .A2(new_n632), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT34), .B(G104), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND2_X1  g484(.A1(new_n378), .A2(new_n382), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n417), .A2(KEYINPUT20), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n420), .B1(new_n415), .B2(new_n416), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(G475), .B2(new_n424), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n667), .A2(new_n638), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT35), .B(G107), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  INV_X1    g493(.A(new_n595), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT36), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n613), .A2(new_n619), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n629), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n627), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n307), .A2(new_n427), .A3(new_n440), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n494), .A2(new_n662), .A3(new_n666), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT37), .B(G110), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  OAI211_X1 g505(.A(new_n686), .B(new_n438), .C1(new_n637), .C2(new_n305), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n424), .A2(G475), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n433), .B(KEYINPUT101), .Z(new_n695));
  XOR2_X1   g509(.A(KEYINPUT99), .B(G900), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n434), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT100), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n694), .B(new_n699), .C1(new_n672), .C2(new_n673), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n378), .B2(new_n382), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n494), .A3(new_n583), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XNOR2_X1  g517(.A(new_n699), .B(KEYINPUT39), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n494), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT103), .Z(new_n706));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n705), .B(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n301), .A2(new_n306), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT38), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n551), .A2(new_n558), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n509), .A2(new_n511), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n565), .B2(new_n566), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n540), .A2(G472), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n660), .A2(new_n279), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT102), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n686), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n425), .B1(new_n378), .B2(new_n382), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n438), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n712), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n708), .A2(new_n710), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  INV_X1    g541(.A(new_n699), .ZN(new_n728));
  AOI211_X1 g542(.A(new_n425), .B(new_n728), .C1(new_n649), .C2(new_n654), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n693), .A3(new_n583), .A4(new_n494), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  OAI21_X1  g545(.A(new_n279), .B1(new_n578), .B2(new_n573), .ZN(new_n732));
  INV_X1    g546(.A(new_n572), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT73), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n579), .A2(new_n580), .A3(G472), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n631), .B1(new_n713), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n492), .A2(new_n487), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n482), .A2(new_n469), .B1(new_n490), .B2(new_n447), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n741), .A3(new_n442), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT104), .B1(new_n659), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n647), .A2(new_n641), .A3(new_n648), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT97), .B1(new_n652), .B2(new_n653), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n656), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n655), .A2(new_n640), .A3(new_n656), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n583), .A2(new_n743), .A3(new_n632), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n639), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NOR2_X1   g571(.A1(new_n676), .A2(new_n638), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n738), .A3(new_n743), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  OAI21_X1  g574(.A(new_n438), .B1(new_n637), .B2(new_n305), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n742), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n426), .A2(new_n437), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n583), .A4(new_n686), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  AOI21_X1  g579(.A(new_n439), .B1(new_n298), .B2(new_n300), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n671), .A3(new_n656), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n542), .A2(new_n547), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n559), .A2(new_n567), .A3(new_n569), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n714), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n550), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n631), .A2(new_n661), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n742), .A2(new_n437), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n767), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT105), .B(G122), .Z(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G24));
  NOR3_X1   g590(.A1(new_n722), .A2(new_n771), .A3(new_n661), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n729), .A2(new_n762), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  AOI21_X1  g593(.A(new_n439), .B1(new_n301), .B2(new_n306), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n494), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT106), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n551), .B(new_n782), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n735), .A2(new_n736), .B1(new_n663), .B2(KEYINPUT32), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n631), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n785), .A3(new_n729), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n494), .A3(new_n583), .A4(new_n632), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n729), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT42), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n786), .A2(KEYINPUT42), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G131), .ZN(G33));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n793), .A3(new_n738), .A4(new_n701), .ZN(new_n794));
  INV_X1    g608(.A(new_n701), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT107), .B1(new_n787), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NAND2_X1  g612(.A1(new_n480), .A2(new_n485), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n487), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  INV_X1    g616(.A(new_n488), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT46), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n804), .A2(new_n805), .B1(new_n487), .B2(new_n492), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n442), .A3(new_n704), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT108), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n780), .B(KEYINPUT110), .Z(new_n811));
  AOI21_X1  g625(.A(KEYINPUT109), .B1(new_n655), .B2(new_n425), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n722), .B1(new_n666), .B2(new_n662), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT44), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT44), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n811), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n808), .A2(new_n820), .A3(new_n442), .A4(new_n704), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n810), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G137), .ZN(G39));
  INV_X1    g637(.A(new_n780), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n789), .A2(new_n824), .A3(new_n583), .A4(new_n632), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n808), .A2(KEYINPUT47), .A3(new_n442), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT47), .B1(new_n808), .B2(new_n442), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  NAND2_X1  g644(.A1(new_n428), .A2(new_n240), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n824), .A2(new_n742), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n721), .A2(new_n433), .A3(new_n631), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n656), .A3(new_n655), .ZN(new_n835));
  INV_X1    g649(.A(new_n695), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n813), .A2(new_n836), .A3(new_n814), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n832), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n835), .B1(new_n838), .B2(new_n777), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n837), .A2(new_n772), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n712), .A2(new_n439), .A3(new_n743), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT50), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n772), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n845), .A3(new_n841), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n806), .A2(new_n807), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n443), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n739), .A2(new_n741), .A3(new_n443), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n826), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n844), .A2(new_n811), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(KEYINPUT115), .A3(new_n853), .ZN(new_n857));
  AOI211_X1 g671(.A(KEYINPUT116), .B(KEYINPUT51), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n855), .ZN(new_n860));
  INV_X1    g674(.A(new_n847), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n838), .A2(new_n785), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT48), .ZN(new_n867));
  INV_X1    g681(.A(new_n751), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n431), .B1(new_n834), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n840), .B2(new_n762), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n847), .A2(new_n863), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n854), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n759), .A2(new_n774), .A3(new_n764), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n755), .A2(new_n791), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n780), .A2(new_n494), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n729), .A2(new_n777), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n671), .A2(new_n700), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n583), .A3(new_n686), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n794), .B2(new_n796), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n687), .A2(new_n688), .B1(new_n441), .B2(new_n633), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n301), .A2(new_n306), .A3(new_n440), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n426), .B1(new_n655), .B2(new_n425), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n667), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n882), .A2(new_n887), .A3(KEYINPUT53), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n686), .A2(new_n728), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n767), .A2(new_n494), .A3(new_n721), .A4(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n730), .A3(new_n702), .A4(new_n778), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT52), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n692), .B1(new_n737), .B2(new_n713), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n893), .B(new_n494), .C1(new_n701), .C2(new_n729), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n778), .A4(new_n890), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT113), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT113), .B1(new_n892), .B2(new_n896), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n876), .B(new_n888), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n874), .B1(new_n745), .B2(new_n754), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(new_n791), .A3(new_n887), .A4(new_n882), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n892), .A2(new_n896), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT113), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT113), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n882), .A2(new_n887), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n900), .A3(new_n876), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n903), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n876), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT53), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT54), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n901), .A2(new_n791), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n882), .A2(new_n887), .A3(KEYINPUT53), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT54), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(KEYINPUT114), .A3(new_n904), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n873), .A2(new_n908), .A3(new_n919), .A4(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n831), .B1(new_n865), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n632), .A2(new_n438), .A3(new_n442), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n656), .B1(new_n927), .B2(KEYINPUT111), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(KEYINPUT111), .B2(new_n927), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n739), .A2(new_n741), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(KEYINPUT49), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(KEYINPUT49), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT112), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n721), .B1(new_n649), .B2(new_n654), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n931), .A2(new_n712), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n935), .ZN(G75));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n899), .A2(new_n904), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(G902), .ZN(new_n939));
  INV_X1    g753(.A(G210), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n239), .A2(new_n276), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n274), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT55), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n944), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n937), .B(new_n946), .C1(new_n939), .C2(new_n940), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n240), .A2(G952), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT117), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G51));
  XOR2_X1   g766(.A(new_n802), .B(KEYINPUT120), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n939), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n803), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT119), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n899), .A2(new_n904), .A3(new_n957), .A4(new_n905), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n916), .A2(new_n900), .B1(new_n912), .B2(new_n922), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n905), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n923), .B2(new_n904), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n740), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT121), .B1(new_n964), .B2(new_n948), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT121), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n906), .A2(KEYINPUT119), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n967), .B(new_n958), .C1(new_n905), .C2(new_n959), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n740), .B1(new_n968), .B2(new_n956), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n966), .B(new_n949), .C1(new_n969), .C2(new_n954), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n965), .A2(new_n970), .ZN(G54));
  AND4_X1   g785(.A1(KEYINPUT58), .A2(new_n938), .A3(G475), .A4(G902), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n949), .B1(new_n972), .B2(new_n415), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n415), .B2(new_n972), .ZN(G60));
  NAND2_X1  g788(.A1(new_n644), .A2(new_n646), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n919), .A2(new_n908), .A3(new_n924), .ZN(new_n976));
  NAND2_X1  g790(.A1(G478), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT59), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n975), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n968), .A2(new_n975), .A3(new_n978), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n948), .ZN(G63));
  XNOR2_X1  g795(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n982));
  OR3_X1    g796(.A1(new_n309), .A2(new_n279), .A3(KEYINPUT60), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT60), .B1(new_n309), .B2(new_n279), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n938), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n949), .B1(new_n985), .B2(new_n628), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n684), .A2(new_n938), .A3(new_n983), .A4(new_n984), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n992), .B(new_n982), .C1(new_n986), .C2(new_n987), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(G66));
  INV_X1    g808(.A(G224), .ZN(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n435), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n901), .A2(new_n887), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n998), .B2(G953), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n942), .B1(G898), .B2(new_n240), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT124), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n999), .B(new_n1001), .ZN(G69));
  AOI21_X1  g816(.A(new_n240), .B1(G227), .B2(G900), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n810), .A2(new_n767), .A3(new_n785), .A4(new_n821), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n894), .A2(new_n778), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n791), .A2(new_n1005), .A3(new_n797), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1004), .A2(new_n822), .A3(new_n829), .A4(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n545), .B1(new_n533), .B2(new_n524), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT125), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(new_n409), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1007), .A2(new_n240), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n738), .A2(new_n780), .ZN(new_n1012));
  INV_X1    g826(.A(new_n885), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(KEYINPUT126), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n706), .B(new_n1014), .C1(KEYINPUT126), .C2(new_n1013), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n726), .A2(KEYINPUT62), .A3(new_n1005), .ZN(new_n1016));
  AOI21_X1  g830(.A(KEYINPUT62), .B1(new_n726), .B2(new_n1005), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n822), .A2(new_n829), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1020), .A2(G953), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1011), .B1(new_n1021), .B2(new_n1010), .ZN(new_n1022));
  INV_X1    g836(.A(G900), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1003), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1003), .B2(new_n1022), .ZN(G72));
  NOR2_X1   g839(.A1(new_n1007), .A2(new_n997), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n717), .B(KEYINPUT63), .Z(new_n1027));
  OAI211_X1 g841(.A(new_n538), .B(new_n546), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n546), .A2(new_n538), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1018), .A2(new_n1019), .A3(new_n997), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n538), .B1(new_n555), .B2(new_n527), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1027), .B1(new_n1032), .B2(new_n540), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n948), .B1(new_n918), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1028), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(KEYINPUT127), .ZN(new_n1036));
  INV_X1    g850(.A(KEYINPUT127), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1028), .A2(new_n1031), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1036), .A2(new_n1038), .ZN(G57));
endmodule


