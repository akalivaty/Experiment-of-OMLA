

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751;

  XNOR2_X1 U379 ( .A(n472), .B(n410), .ZN(n726) );
  XNOR2_X1 U380 ( .A(n449), .B(G128), .ZN(n484) );
  XNOR2_X1 U381 ( .A(n460), .B(n459), .ZN(n461) );
  NOR2_X1 U382 ( .A1(n551), .A2(n603), .ZN(n552) );
  NOR2_X1 U383 ( .A1(n620), .A2(n619), .ZN(n653) );
  XNOR2_X1 U384 ( .A(n484), .B(n448), .ZN(n732) );
  XNOR2_X1 U385 ( .A(n431), .B(n582), .ZN(n589) );
  NOR2_X1 U386 ( .A1(n570), .A2(n562), .ZN(n637) );
  AND2_X2 U387 ( .A1(n436), .A2(n358), .ZN(n733) );
  XNOR2_X2 U388 ( .A(n377), .B(n435), .ZN(n436) );
  XNOR2_X2 U389 ( .A(n599), .B(KEYINPUT35), .ZN(n607) );
  NOR2_X2 U390 ( .A1(n749), .A2(n750), .ZN(n401) );
  XNOR2_X2 U391 ( .A(n397), .B(n396), .ZN(n749) );
  XNOR2_X2 U392 ( .A(n505), .B(G125), .ZN(n472) );
  XNOR2_X1 U393 ( .A(n548), .B(KEYINPUT79), .ZN(n561) );
  XNOR2_X1 U394 ( .A(n574), .B(n437), .ZN(n603) );
  INV_X4 U395 ( .A(G146), .ZN(n505) );
  AND2_X1 U396 ( .A1(n375), .A2(n373), .ZN(n372) );
  NOR2_X1 U397 ( .A1(n693), .A2(G953), .ZN(n399) );
  AND2_X2 U398 ( .A1(n622), .A2(n621), .ZN(n707) );
  NAND2_X1 U399 ( .A1(n380), .A2(n379), .ZN(n610) );
  AND2_X1 U400 ( .A1(n381), .A2(n382), .ZN(n380) );
  XNOR2_X1 U401 ( .A(n441), .B(n440), .ZN(n747) );
  NOR2_X1 U402 ( .A1(n391), .A2(n585), .ZN(n629) );
  NAND2_X1 U403 ( .A1(n561), .A2(n668), .ZN(n549) );
  AND2_X1 U404 ( .A1(n389), .A2(n427), .ZN(n605) );
  OR2_X1 U405 ( .A1(n584), .A2(n595), .ZN(n585) );
  NOR2_X1 U406 ( .A1(n603), .A2(n593), .ZN(n594) );
  NAND2_X1 U407 ( .A1(n378), .A2(n580), .ZN(n431) );
  XNOR2_X1 U408 ( .A(n556), .B(KEYINPUT19), .ZN(n378) );
  NAND2_X1 U409 ( .A1(n550), .A2(n669), .ZN(n556) );
  XNOR2_X1 U410 ( .A(n456), .B(G107), .ZN(n718) );
  XNOR2_X1 U411 ( .A(G116), .B(KEYINPUT73), .ZN(n458) );
  XNOR2_X1 U412 ( .A(G104), .B(G110), .ZN(n456) );
  INV_X1 U413 ( .A(G134), .ZN(n448) );
  XNOR2_X1 U414 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U415 ( .A(KEYINPUT70), .ZN(n403) );
  XNOR2_X1 U416 ( .A(G137), .B(KEYINPUT69), .ZN(n533) );
  INV_X1 U417 ( .A(G143), .ZN(n449) );
  XNOR2_X1 U418 ( .A(n552), .B(KEYINPUT102), .ZN(n426) );
  INV_X1 U419 ( .A(G472), .ZN(n438) );
  NAND2_X1 U420 ( .A1(n707), .A2(n413), .ZN(n376) );
  NOR2_X1 U421 ( .A1(n627), .A2(n414), .ZN(n413) );
  INV_X1 U422 ( .A(G475), .ZN(n414) );
  XNOR2_X1 U423 ( .A(n493), .B(G478), .ZN(n559) );
  NOR2_X1 U424 ( .A1(n633), .A2(n748), .ZN(n608) );
  XNOR2_X1 U425 ( .A(G101), .B(n728), .ZN(n496) );
  XNOR2_X1 U426 ( .A(n607), .B(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U427 ( .A(n383), .B(KEYINPUT99), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n432), .B(n496), .ZN(n530) );
  INV_X1 U429 ( .A(n718), .ZN(n432) );
  INV_X1 U430 ( .A(KEYINPUT48), .ZN(n435) );
  XNOR2_X1 U431 ( .A(n468), .B(KEYINPUT87), .ZN(n469) );
  XNOR2_X1 U432 ( .A(n539), .B(G469), .ZN(n450) );
  XNOR2_X1 U433 ( .A(KEYINPUT16), .B(G122), .ZN(n463) );
  XOR2_X1 U434 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n464) );
  XNOR2_X1 U435 ( .A(n513), .B(n409), .ZN(n408) );
  XNOR2_X1 U436 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n513) );
  XNOR2_X1 U437 ( .A(KEYINPUT89), .B(KEYINPUT75), .ZN(n409) );
  XNOR2_X1 U438 ( .A(n407), .B(G140), .ZN(n406) );
  INV_X1 U439 ( .A(G110), .ZN(n407) );
  XNOR2_X1 U440 ( .A(G119), .B(G128), .ZN(n515) );
  INV_X1 U441 ( .A(KEYINPUT10), .ZN(n410) );
  XNOR2_X1 U442 ( .A(G107), .B(KEYINPUT9), .ZN(n485) );
  XOR2_X1 U443 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n486) );
  XNOR2_X1 U444 ( .A(n732), .B(n362), .ZN(n395) );
  NOR2_X1 U445 ( .A1(n418), .A2(n419), .ZN(n443) );
  NOR2_X1 U446 ( .A1(n426), .A2(n553), .ZN(n419) );
  NAND2_X1 U447 ( .A1(n422), .A2(n420), .ZN(n418) );
  AND2_X1 U448 ( .A1(n421), .A2(n424), .ZN(n420) );
  INV_X1 U449 ( .A(KEYINPUT6), .ZN(n437) );
  XNOR2_X1 U450 ( .A(n523), .B(n360), .ZN(n434) );
  NOR2_X1 U451 ( .A1(n709), .A2(G902), .ZN(n523) );
  XNOR2_X1 U452 ( .A(n590), .B(n390), .ZN(n389) );
  INV_X1 U453 ( .A(KEYINPUT22), .ZN(n390) );
  NOR2_X1 U454 ( .A1(n707), .A2(n417), .ZN(n415) );
  NAND2_X1 U455 ( .A1(n374), .A2(n367), .ZN(n373) );
  NAND2_X1 U456 ( .A1(n376), .A2(n411), .ZN(n374) );
  NOR2_X1 U457 ( .A1(n370), .A2(n367), .ZN(n369) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n564) );
  INV_X1 U459 ( .A(KEYINPUT47), .ZN(n392) );
  NOR2_X1 U460 ( .A1(n639), .A2(n673), .ZN(n393) );
  XOR2_X1 U461 ( .A(G104), .B(G122), .Z(n477) );
  XNOR2_X1 U462 ( .A(G113), .B(G143), .ZN(n476) );
  XNOR2_X1 U463 ( .A(n452), .B(G140), .ZN(n534) );
  INV_X1 U464 ( .A(G131), .ZN(n452) );
  OR2_X1 U465 ( .A1(G237), .A2(G902), .ZN(n467) );
  XOR2_X1 U466 ( .A(G137), .B(KEYINPUT93), .Z(n500) );
  XNOR2_X1 U467 ( .A(G131), .B(KEYINPUT5), .ZN(n495) );
  XNOR2_X1 U468 ( .A(n534), .B(n533), .ZN(n727) );
  XNOR2_X1 U469 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  XNOR2_X1 U470 ( .A(n732), .B(n505), .ZN(n531) );
  XNOR2_X1 U471 ( .A(n727), .B(n451), .ZN(n454) );
  INV_X1 U472 ( .A(KEYINPUT81), .ZN(n451) );
  NAND2_X1 U473 ( .A1(G234), .A2(G237), .ZN(n507) );
  XOR2_X1 U474 ( .A(n471), .B(n550), .Z(n668) );
  OR2_X1 U475 ( .A1(n425), .A2(n553), .ZN(n421) );
  INV_X1 U476 ( .A(n556), .ZN(n424) );
  NAND2_X1 U477 ( .A1(n426), .A2(n423), .ZN(n422) );
  NAND2_X1 U478 ( .A1(n657), .A2(n656), .ZN(n593) );
  NOR2_X1 U479 ( .A1(n542), .A2(n584), .ZN(n543) );
  NOR2_X1 U480 ( .A1(n542), .A2(n527), .ZN(n528) );
  XNOR2_X1 U481 ( .A(n483), .B(n482), .ZN(n560) );
  AND2_X1 U482 ( .A1(n434), .A2(n428), .ZN(n656) );
  INV_X1 U483 ( .A(n587), .ZN(n428) );
  NAND2_X1 U484 ( .A1(n359), .A2(n385), .ZN(n379) );
  NOR2_X1 U485 ( .A1(n412), .A2(n711), .ZN(n411) );
  NOR2_X1 U486 ( .A1(n417), .A2(G475), .ZN(n412) );
  XNOR2_X1 U487 ( .A(n387), .B(n530), .ZN(n386) );
  XNOR2_X1 U488 ( .A(n455), .B(n388), .ZN(n387) );
  XNOR2_X1 U489 ( .A(n484), .B(n466), .ZN(n388) );
  XNOR2_X1 U490 ( .A(n519), .B(n518), .ZN(n709) );
  XNOR2_X1 U491 ( .A(n726), .B(n405), .ZN(n519) );
  XNOR2_X1 U492 ( .A(n408), .B(n406), .ZN(n405) );
  XNOR2_X1 U493 ( .A(n488), .B(n395), .ZN(n492) );
  XNOR2_X1 U494 ( .A(n541), .B(KEYINPUT42), .ZN(n750) );
  INV_X1 U495 ( .A(KEYINPUT40), .ZN(n396) );
  INV_X1 U496 ( .A(KEYINPUT107), .ZN(n440) );
  NAND2_X1 U497 ( .A1(n442), .A2(n657), .ZN(n441) );
  NAND2_X1 U498 ( .A1(n603), .A2(n434), .ZN(n433) );
  NAND2_X1 U499 ( .A1(n371), .A2(n363), .ZN(n368) );
  INV_X1 U500 ( .A(n415), .ZN(n371) );
  INV_X1 U501 ( .A(KEYINPUT56), .ZN(n444) );
  AND2_X1 U502 ( .A1(n744), .A2(n616), .ZN(n358) );
  AND2_X1 U503 ( .A1(n608), .A2(n600), .ZN(n359) );
  INV_X1 U504 ( .A(n640), .ZN(n425) );
  XOR2_X1 U505 ( .A(n522), .B(n521), .Z(n360) );
  AND2_X1 U506 ( .A1(n426), .A2(n425), .ZN(n361) );
  XOR2_X1 U507 ( .A(G116), .B(G122), .Z(n362) );
  AND2_X1 U508 ( .A1(n376), .A2(n369), .ZN(n363) );
  NOR2_X1 U509 ( .A1(n433), .A2(n657), .ZN(n364) );
  XNOR2_X1 U510 ( .A(n386), .B(n719), .ZN(n694) );
  XOR2_X1 U511 ( .A(n696), .B(n695), .Z(n365) );
  XOR2_X1 U512 ( .A(n624), .B(KEYINPUT62), .Z(n366) );
  INV_X1 U513 ( .A(n627), .ZN(n417) );
  XOR2_X1 U514 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n367) );
  NOR2_X1 U515 ( .A1(G952), .A2(n735), .ZN(n711) );
  INV_X1 U516 ( .A(n711), .ZN(n416) );
  NAND2_X1 U517 ( .A1(n372), .A2(n368), .ZN(G60) );
  INV_X1 U518 ( .A(n411), .ZN(n370) );
  NAND2_X1 U519 ( .A1(n415), .A2(n367), .ZN(n375) );
  NAND2_X1 U520 ( .A1(n400), .A2(n402), .ZN(n377) );
  NAND2_X1 U521 ( .A1(n558), .A2(n378), .ZN(n639) );
  OR2_X1 U522 ( .A1(n592), .A2(n751), .ZN(n383) );
  NAND2_X1 U523 ( .A1(n384), .A2(KEYINPUT44), .ZN(n381) );
  NAND2_X1 U524 ( .A1(n609), .A2(n608), .ZN(n384) );
  NAND2_X1 U525 ( .A1(n694), .A2(n611), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n502), .B(n465), .ZN(n719) );
  AND2_X1 U527 ( .A1(n389), .A2(n364), .ZN(n591) );
  NAND2_X1 U528 ( .A1(n436), .A2(n744), .ZN(n620) );
  XNOR2_X1 U529 ( .A(n447), .B(n365), .ZN(n446) );
  OR2_X1 U530 ( .A1(n615), .A2(n614), .ZN(n622) );
  NOR2_X1 U531 ( .A1(n601), .A2(n551), .ZN(n529) );
  NAND2_X1 U532 ( .A1(n446), .A2(n416), .ZN(n445) );
  NAND2_X1 U533 ( .A1(n707), .A2(G210), .ZN(n447) );
  INV_X1 U534 ( .A(n574), .ZN(n663) );
  XNOR2_X2 U535 ( .A(n439), .B(n438), .ZN(n574) );
  NOR2_X1 U536 ( .A1(n697), .A2(G902), .ZN(n538) );
  BUF_X1 U537 ( .A(n663), .Z(n391) );
  NAND2_X1 U538 ( .A1(n394), .A2(n540), .ZN(n557) );
  XNOR2_X1 U539 ( .A(n529), .B(KEYINPUT28), .ZN(n394) );
  XNOR2_X1 U540 ( .A(n443), .B(KEYINPUT36), .ZN(n442) );
  NAND2_X1 U541 ( .A1(n573), .A2(n425), .ZN(n397) );
  NAND2_X1 U542 ( .A1(n398), .A2(n547), .ZN(n548) );
  XNOR2_X1 U543 ( .A(n546), .B(n545), .ZN(n398) );
  XNOR2_X1 U544 ( .A(n399), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U545 ( .A(n401), .B(KEYINPUT46), .ZN(n400) );
  XNOR2_X1 U546 ( .A(n503), .B(n504), .ZN(n506) );
  NAND2_X1 U547 ( .A1(n544), .A2(n669), .ZN(n546) );
  XNOR2_X2 U548 ( .A(n663), .B(KEYINPUT100), .ZN(n544) );
  XNOR2_X1 U549 ( .A(n445), .B(n444), .ZN(G51) );
  NAND2_X1 U550 ( .A1(n565), .A2(n747), .ZN(n404) );
  AND2_X1 U551 ( .A1(n425), .A2(n553), .ZN(n423) );
  NAND2_X1 U552 ( .A1(n427), .A2(n654), .ZN(n527) );
  INV_X1 U553 ( .A(n434), .ZN(n427) );
  OR2_X2 U554 ( .A1(n623), .A2(G902), .ZN(n439) );
  XNOR2_X2 U555 ( .A(n549), .B(KEYINPUT39), .ZN(n573) );
  XNOR2_X1 U556 ( .A(n429), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U557 ( .A1(n430), .A2(n416), .ZN(n429) );
  XNOR2_X1 U558 ( .A(n625), .B(n366), .ZN(n430) );
  XNOR2_X2 U559 ( .A(n554), .B(KEYINPUT1), .ZN(n657) );
  XNOR2_X2 U560 ( .A(n538), .B(n450), .ZN(n554) );
  XNOR2_X1 U561 ( .A(n532), .B(n531), .ZN(n537) );
  XNOR2_X2 U562 ( .A(G119), .B(KEYINPUT3), .ZN(n460) );
  INV_X1 U563 ( .A(n530), .ZN(n532) );
  XOR2_X1 U564 ( .A(n477), .B(n476), .Z(n453) );
  XOR2_X1 U565 ( .A(n457), .B(n472), .Z(n455) );
  INV_X1 U566 ( .A(KEYINPUT74), .ZN(n459) );
  INV_X1 U567 ( .A(KEYINPUT30), .ZN(n545) );
  XNOR2_X1 U568 ( .A(n478), .B(n453), .ZN(n479) );
  XNOR2_X1 U569 ( .A(n481), .B(G475), .ZN(n482) );
  XNOR2_X1 U570 ( .A(n480), .B(n479), .ZN(n626) );
  INV_X1 U571 ( .A(n657), .ZN(n567) );
  XNOR2_X1 U572 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U573 ( .A(n544), .ZN(n601) );
  NAND2_X1 U574 ( .A1(G214), .A2(n467), .ZN(n669) );
  XNOR2_X1 U575 ( .A(KEYINPUT38), .B(KEYINPUT78), .ZN(n471) );
  XNOR2_X2 U576 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n728) );
  INV_X2 U577 ( .A(G953), .ZN(n735) );
  AND2_X1 U578 ( .A1(G224), .A2(n735), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n458), .B(G113), .ZN(n462) );
  XNOR2_X2 U580 ( .A(n462), .B(n461), .ZN(n502) );
  XNOR2_X1 U581 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U582 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n466) );
  NAND2_X1 U583 ( .A1(G210), .A2(n467), .ZN(n468) );
  XNOR2_X2 U584 ( .A(n470), .B(n469), .ZN(n550) );
  NAND2_X1 U585 ( .A1(n669), .A2(n668), .ZN(n672) );
  XNOR2_X1 U586 ( .A(n534), .B(n726), .ZN(n480) );
  XOR2_X1 U587 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n474) );
  NOR2_X1 U588 ( .A1(G953), .A2(G237), .ZN(n498) );
  NAND2_X1 U589 ( .A1(G214), .A2(n498), .ZN(n473) );
  XNOR2_X1 U590 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U591 ( .A(n475), .B(KEYINPUT94), .Z(n478) );
  NOR2_X1 U592 ( .A1(G902), .A2(n626), .ZN(n483) );
  XNOR2_X1 U593 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U595 ( .A(n487), .B(KEYINPUT96), .Z(n488) );
  XOR2_X1 U596 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n490) );
  NAND2_X1 U597 ( .A1(G234), .A2(n735), .ZN(n489) );
  XNOR2_X1 U598 ( .A(n490), .B(n489), .ZN(n514) );
  NAND2_X1 U599 ( .A1(G217), .A2(n514), .ZN(n491) );
  XNOR2_X1 U600 ( .A(n492), .B(n491), .ZN(n703) );
  NOR2_X1 U601 ( .A1(n703), .A2(G902), .ZN(n493) );
  NAND2_X1 U602 ( .A1(n560), .A2(n559), .ZN(n671) );
  NOR2_X1 U603 ( .A1(n672), .A2(n671), .ZN(n494) );
  XNOR2_X1 U604 ( .A(n494), .B(KEYINPUT41), .ZN(n685) );
  XNOR2_X1 U605 ( .A(n495), .B(KEYINPUT92), .ZN(n497) );
  XOR2_X1 U606 ( .A(n497), .B(n496), .Z(n504) );
  NAND2_X1 U607 ( .A1(n498), .A2(G210), .ZN(n499) );
  XNOR2_X1 U608 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U609 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U610 ( .A(n506), .B(n531), .ZN(n623) );
  XNOR2_X1 U611 ( .A(n507), .B(KEYINPUT14), .ZN(n509) );
  NAND2_X1 U612 ( .A1(G952), .A2(n509), .ZN(n508) );
  XNOR2_X1 U613 ( .A(KEYINPUT88), .B(n508), .ZN(n683) );
  NOR2_X1 U614 ( .A1(G953), .A2(n683), .ZN(n577) );
  NAND2_X1 U615 ( .A1(G902), .A2(n509), .ZN(n575) );
  NOR2_X1 U616 ( .A1(G900), .A2(n575), .ZN(n510) );
  NAND2_X1 U617 ( .A1(G953), .A2(n510), .ZN(n511) );
  XNOR2_X1 U618 ( .A(KEYINPUT101), .B(n511), .ZN(n512) );
  NOR2_X1 U619 ( .A1(n577), .A2(n512), .ZN(n542) );
  AND2_X1 U620 ( .A1(G221), .A2(n514), .ZN(n517) );
  XOR2_X1 U621 ( .A(n515), .B(n533), .Z(n516) );
  NAND2_X1 U622 ( .A1(n611), .A2(G234), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n520), .B(KEYINPUT20), .ZN(n524) );
  NAND2_X1 U624 ( .A1(G217), .A2(n524), .ZN(n522) );
  INV_X1 U625 ( .A(KEYINPUT25), .ZN(n521) );
  XOR2_X1 U626 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n526) );
  NAND2_X1 U627 ( .A1(n524), .A2(G221), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n526), .B(n525), .ZN(n654) );
  XNOR2_X1 U629 ( .A(n528), .B(KEYINPUT71), .ZN(n551) );
  INV_X1 U630 ( .A(KEYINPUT72), .ZN(n539) );
  NAND2_X1 U631 ( .A1(G227), .A2(n735), .ZN(n535) );
  XNOR2_X1 U632 ( .A(n454), .B(n535), .ZN(n536) );
  XNOR2_X1 U633 ( .A(n537), .B(n536), .ZN(n697) );
  XOR2_X1 U634 ( .A(n554), .B(KEYINPUT105), .Z(n540) );
  NOR2_X1 U635 ( .A1(n685), .A2(n557), .ZN(n541) );
  INV_X1 U636 ( .A(n560), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n555), .A2(n559), .ZN(n640) );
  XNOR2_X1 U638 ( .A(n654), .B(KEYINPUT91), .ZN(n587) );
  NAND2_X1 U639 ( .A1(n656), .A2(n554), .ZN(n584) );
  XNOR2_X1 U640 ( .A(n543), .B(KEYINPUT80), .ZN(n547) );
  INV_X1 U641 ( .A(KEYINPUT106), .ZN(n553) );
  NOR2_X1 U642 ( .A1(n555), .A2(n559), .ZN(n644) );
  NOR2_X1 U643 ( .A1(n425), .A2(n644), .ZN(n673) );
  INV_X1 U644 ( .A(n557), .ZN(n558) );
  INV_X1 U645 ( .A(n550), .ZN(n570) );
  NOR2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n597) );
  NAND2_X1 U647 ( .A1(n561), .A2(n597), .ZN(n562) );
  XNOR2_X1 U648 ( .A(n637), .B(KEYINPUT84), .ZN(n563) );
  NOR2_X1 U649 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U650 ( .A1(n361), .A2(n669), .ZN(n566) );
  XNOR2_X1 U651 ( .A(n566), .B(KEYINPUT103), .ZN(n568) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n569), .B(KEYINPUT43), .ZN(n571) );
  NAND2_X1 U654 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U655 ( .A(KEYINPUT104), .B(n572), .ZN(n744) );
  NAND2_X1 U656 ( .A1(n644), .A2(n573), .ZN(n616) );
  INV_X1 U657 ( .A(n616), .ZN(n649) );
  NOR2_X1 U658 ( .A1(n574), .A2(n593), .ZN(n665) );
  NOR2_X1 U659 ( .A1(G898), .A2(n735), .ZN(n722) );
  INV_X1 U660 ( .A(n575), .ZN(n576) );
  NAND2_X1 U661 ( .A1(n722), .A2(n576), .ZN(n579) );
  INV_X1 U662 ( .A(n577), .ZN(n578) );
  NAND2_X1 U663 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U664 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n581) );
  XOR2_X1 U665 ( .A(KEYINPUT66), .B(n581), .Z(n582) );
  INV_X1 U666 ( .A(n589), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n665), .A2(n589), .ZN(n583) );
  XNOR2_X1 U668 ( .A(n583), .B(KEYINPUT31), .ZN(n645) );
  NOR2_X1 U669 ( .A1(n645), .A2(n629), .ZN(n586) );
  NOR2_X1 U670 ( .A1(n673), .A2(n586), .ZN(n592) );
  NOR2_X1 U671 ( .A1(n587), .A2(n671), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U673 ( .A(KEYINPUT98), .B(n591), .ZN(n751) );
  XNOR2_X1 U674 ( .A(KEYINPUT33), .B(n594), .ZN(n684) );
  NOR2_X1 U675 ( .A1(n595), .A2(n684), .ZN(n596) );
  XNOR2_X1 U676 ( .A(n596), .B(KEYINPUT34), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U678 ( .A(KEYINPUT44), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n605), .A2(n601), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n657), .A2(n602), .ZN(n633) );
  AND2_X1 U681 ( .A1(n603), .A2(n657), .ZN(n604) );
  AND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(KEYINPUT32), .ZN(n748) );
  NOR2_X1 U684 ( .A1(n607), .A2(KEYINPUT67), .ZN(n609) );
  XNOR2_X2 U685 ( .A(n610), .B(KEYINPUT45), .ZN(n715) );
  NAND2_X1 U686 ( .A1(n733), .A2(n715), .ZN(n650) );
  NOR2_X1 U687 ( .A1(n650), .A2(n611), .ZN(n615) );
  INV_X1 U688 ( .A(n611), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(KEYINPUT65), .ZN(n614) );
  NAND2_X1 U691 ( .A1(KEYINPUT2), .A2(n616), .ZN(n617) );
  XOR2_X1 U692 ( .A(KEYINPUT82), .B(n617), .Z(n618) );
  NAND2_X1 U693 ( .A1(n715), .A2(n618), .ZN(n619) );
  INV_X1 U694 ( .A(n653), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n707), .A2(G472), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n623), .B(KEYINPUT86), .ZN(n624) );
  XOR2_X1 U697 ( .A(n626), .B(KEYINPUT59), .Z(n627) );
  NAND2_X1 U698 ( .A1(n629), .A2(n425), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(G104), .ZN(G6) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n631) );
  NAND2_X1 U701 ( .A1(n629), .A2(n644), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(G107), .B(n632), .ZN(G9) );
  XOR2_X1 U704 ( .A(G110), .B(n633), .Z(G12) );
  INV_X1 U705 ( .A(n644), .ZN(n634) );
  NOR2_X1 U706 ( .A1(n634), .A2(n639), .ZN(n636) );
  XNOR2_X1 U707 ( .A(G128), .B(KEYINPUT29), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G30) );
  XOR2_X1 U709 ( .A(G143), .B(n637), .Z(n638) );
  XNOR2_X1 U710 ( .A(KEYINPUT108), .B(n638), .ZN(G45) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U712 ( .A(G146), .B(KEYINPUT109), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G48) );
  NAND2_X1 U714 ( .A1(n645), .A2(n425), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(G113), .ZN(G15) );
  XOR2_X1 U716 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n647) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(G116), .B(n648), .ZN(G18) );
  XOR2_X1 U720 ( .A(G134), .B(n649), .Z(G36) );
  INV_X1 U721 ( .A(n650), .ZN(n651) );
  NOR2_X1 U722 ( .A1(KEYINPUT2), .A2(n651), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n691) );
  NOR2_X1 U724 ( .A1(n654), .A2(n434), .ZN(n655) );
  XNOR2_X1 U725 ( .A(KEYINPUT49), .B(n655), .ZN(n661) );
  XNOR2_X1 U726 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n391), .A2(n662), .ZN(n664) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n666), .Z(n667) );
  NOR2_X1 U733 ( .A1(n685), .A2(n667), .ZN(n680) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n676) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U737 ( .A(n674), .B(KEYINPUT114), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n677), .A2(n684), .ZN(n678) );
  XOR2_X1 U740 ( .A(KEYINPUT115), .B(n678), .Z(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U742 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n688) );
  NOR2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n686), .B(KEYINPUT116), .ZN(n687) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U747 ( .A(n689), .B(KEYINPUT117), .ZN(n690) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U749 ( .A(KEYINPUT118), .B(n692), .Z(n693) );
  XOR2_X1 U750 ( .A(KEYINPUT83), .B(KEYINPUT55), .Z(n696) );
  XNOR2_X1 U751 ( .A(n694), .B(KEYINPUT54), .ZN(n695) );
  XNOR2_X1 U752 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n697), .B(KEYINPUT57), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U755 ( .A1(n707), .A2(G469), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n711), .A2(n702), .ZN(G54) );
  XOR2_X1 U758 ( .A(n703), .B(KEYINPUT121), .Z(n705) );
  NAND2_X1 U759 ( .A1(n707), .A2(G478), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U761 ( .A1(n711), .A2(n706), .ZN(G63) );
  NAND2_X1 U762 ( .A1(G217), .A2(n707), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(G66) );
  NAND2_X1 U765 ( .A1(G224), .A2(G953), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT122), .ZN(n713) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U768 ( .A1(G898), .A2(n714), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n715), .A2(n735), .ZN(n716) );
  NAND2_X1 U770 ( .A1(n717), .A2(n716), .ZN(n724) );
  XNOR2_X1 U771 ( .A(n718), .B(G101), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U774 ( .A(n724), .B(n723), .Z(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT123), .B(n725), .ZN(G69) );
  XNOR2_X1 U776 ( .A(n726), .B(KEYINPUT124), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U778 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n732), .B(n731), .ZN(n738) );
  XOR2_X1 U780 ( .A(n733), .B(KEYINPUT125), .Z(n734) );
  XNOR2_X1 U781 ( .A(n738), .B(n734), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n736), .A2(n735), .ZN(n743) );
  XOR2_X1 U783 ( .A(G227), .B(KEYINPUT126), .Z(n737) );
  XNOR2_X1 U784 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(G953), .ZN(n741) );
  XOR2_X1 U787 ( .A(KEYINPUT127), .B(n741), .Z(n742) );
  NAND2_X1 U788 ( .A1(n743), .A2(n742), .ZN(G72) );
  XNOR2_X1 U789 ( .A(G140), .B(n744), .ZN(n745) );
  XNOR2_X1 U790 ( .A(n745), .B(KEYINPUT112), .ZN(G42) );
  XOR2_X1 U791 ( .A(n607), .B(G122), .Z(G24) );
  XOR2_X1 U792 ( .A(G125), .B(KEYINPUT37), .Z(n746) );
  XNOR2_X1 U793 ( .A(n747), .B(n746), .ZN(G27) );
  XOR2_X1 U794 ( .A(G119), .B(n748), .Z(G21) );
  XOR2_X1 U795 ( .A(n749), .B(G131), .Z(G33) );
  XOR2_X1 U796 ( .A(G137), .B(n750), .Z(G39) );
  XOR2_X1 U797 ( .A(G101), .B(n751), .Z(G3) );
endmodule

