

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U323 ( .A1(n533), .A2(n457), .ZN(n422) );
  AND2_X1 U324 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U325 ( .A(n343), .B(n291), .ZN(n344) );
  INV_X1 U326 ( .A(KEYINPUT54), .ZN(n421) );
  XNOR2_X1 U327 ( .A(n345), .B(n344), .ZN(n350) );
  XNOR2_X1 U328 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U329 ( .A(n440), .B(KEYINPUT55), .ZN(n453) );
  XNOR2_X1 U330 ( .A(n352), .B(n351), .ZN(n576) );
  XNOR2_X1 U331 ( .A(KEYINPUT41), .B(n576), .ZN(n562) );
  XOR2_X1 U332 ( .A(n467), .B(KEYINPUT28), .Z(n536) );
  XNOR2_X1 U333 ( .A(n454), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U334 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(G43GAT), .B(G134GAT), .Z(n441) );
  XNOR2_X1 U336 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n292), .B(KEYINPUT71), .ZN(n359) );
  XNOR2_X1 U338 ( .A(n441), .B(n359), .ZN(n294) );
  AND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U341 ( .A(KEYINPUT66), .B(KEYINPUT64), .Z(n296) );
  XNOR2_X1 U342 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U345 ( .A(G92GAT), .B(G85GAT), .Z(n300) );
  XNOR2_X1 U346 ( .A(G29GAT), .B(G162GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U349 ( .A(KEYINPUT76), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U350 ( .A(G50GAT), .B(G190GAT), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U353 ( .A(KEYINPUT73), .B(G106GAT), .Z(n308) );
  XNOR2_X1 U354 ( .A(G36GAT), .B(G99GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n310) );
  XNOR2_X1 U357 ( .A(KEYINPUT10), .B(KEYINPUT77), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U360 ( .A(n314), .B(n313), .Z(n559) );
  XOR2_X1 U361 ( .A(G120GAT), .B(G127GAT), .Z(n316) );
  XNOR2_X1 U362 ( .A(KEYINPUT0), .B(KEYINPUT85), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(G113GAT), .B(n317), .Z(n449) );
  XOR2_X1 U365 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n319) );
  XNOR2_X1 U366 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U368 ( .A(n320), .B(G148GAT), .Z(n322) );
  XOR2_X1 U369 ( .A(G29GAT), .B(G1GAT), .Z(n362) );
  XNOR2_X1 U370 ( .A(n362), .B(G134GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U372 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n324) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U375 ( .A(n326), .B(n325), .Z(n331) );
  XOR2_X1 U376 ( .A(G155GAT), .B(G162GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U379 ( .A(G141GAT), .B(n329), .ZN(n438) );
  XOR2_X1 U380 ( .A(G85GAT), .B(G57GAT), .Z(n337) );
  XOR2_X1 U381 ( .A(n438), .B(n337), .Z(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U383 ( .A(n449), .B(n332), .Z(n471) );
  XOR2_X1 U384 ( .A(KEYINPUT96), .B(n471), .Z(n522) );
  INV_X1 U385 ( .A(n559), .ZN(n395) );
  XOR2_X1 U386 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n334) );
  XNOR2_X1 U387 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n352) );
  XNOR2_X1 U389 ( .A(G92GAT), .B(G64GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n335), .B(G204GAT), .ZN(n403) );
  INV_X1 U391 ( .A(n337), .ZN(n336) );
  NAND2_X1 U392 ( .A1(n403), .A2(n336), .ZN(n340) );
  INV_X1 U393 ( .A(n403), .ZN(n338) );
  NAND2_X1 U394 ( .A1(n338), .A2(n337), .ZN(n339) );
  NAND2_X1 U395 ( .A1(n340), .A2(n339), .ZN(n345) );
  XOR2_X1 U396 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n342) );
  XNOR2_X1 U397 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G71GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n346), .B(G176GAT), .ZN(n442) );
  XOR2_X1 U401 ( .A(KEYINPUT72), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U402 ( .A(G148GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n431) );
  XNOR2_X1 U404 ( .A(n442), .B(n431), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U406 ( .A(KEYINPUT29), .B(G113GAT), .Z(n354) );
  XNOR2_X1 U407 ( .A(G197GAT), .B(G141GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U409 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n356) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(KEYINPUT68), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n358), .B(n357), .Z(n369) );
  XOR2_X1 U413 ( .A(n359), .B(KEYINPUT69), .Z(n361) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G43GAT), .Z(n364) );
  XOR2_X1 U417 ( .A(G50GAT), .B(G22GAT), .Z(n430) );
  XNOR2_X1 U418 ( .A(n362), .B(n430), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U421 ( .A(G36GAT), .B(G8GAT), .Z(n410) );
  XOR2_X1 U422 ( .A(n367), .B(n410), .Z(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n507) );
  INV_X1 U424 ( .A(n507), .ZN(n571) );
  NOR2_X1 U425 ( .A1(n562), .A2(n571), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n370), .B(KEYINPUT46), .ZN(n392) );
  XOR2_X1 U427 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n372) );
  XNOR2_X1 U428 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n391) );
  XOR2_X1 U430 ( .A(G211GAT), .B(G64GAT), .Z(n374) );
  XNOR2_X1 U431 ( .A(G1GAT), .B(KEYINPUT13), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U433 ( .A(KEYINPUT82), .B(G78GAT), .Z(n376) );
  XNOR2_X1 U434 ( .A(G127GAT), .B(G155GAT), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U436 ( .A(n378), .B(n377), .Z(n389) );
  XOR2_X1 U437 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n387) );
  XOR2_X1 U440 ( .A(G57GAT), .B(G71GAT), .Z(n382) );
  XNOR2_X1 U441 ( .A(G22GAT), .B(G15GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U443 ( .A(G183GAT), .B(n383), .Z(n385) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n567) );
  INV_X1 U449 ( .A(n567), .ZN(n579) );
  NOR2_X1 U450 ( .A1(n392), .A2(n579), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT118), .B(n393), .Z(n394) );
  NOR2_X1 U452 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n396), .B(KEYINPUT47), .ZN(n401) );
  XNOR2_X1 U454 ( .A(KEYINPUT36), .B(n559), .ZN(n585) );
  OR2_X1 U455 ( .A1(n585), .A2(n567), .ZN(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT45), .B(n397), .ZN(n398) );
  NOR2_X1 U457 ( .A1(n576), .A2(n398), .ZN(n399) );
  NAND2_X1 U458 ( .A1(n399), .A2(n571), .ZN(n400) );
  NAND2_X1 U459 ( .A1(n401), .A2(n400), .ZN(n402) );
  XOR2_X1 U460 ( .A(KEYINPUT48), .B(n402), .Z(n533) );
  XOR2_X1 U461 ( .A(n403), .B(KEYINPUT97), .Z(n405) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n414) );
  XNOR2_X1 U464 ( .A(G218GAT), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n406), .B(KEYINPUT90), .ZN(n407) );
  XOR2_X1 U466 ( .A(n407), .B(KEYINPUT21), .Z(n409) );
  XNOR2_X1 U467 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n435) );
  XOR2_X1 U469 ( .A(n435), .B(KEYINPUT79), .Z(n412) );
  XNOR2_X1 U470 ( .A(n410), .B(G176GAT), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n420) );
  XNOR2_X1 U473 ( .A(KEYINPUT17), .B(G190GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n415), .B(G183GAT), .ZN(n416) );
  XOR2_X1 U475 ( .A(n416), .B(KEYINPUT18), .Z(n418) );
  XNOR2_X1 U476 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n417) );
  XOR2_X1 U477 ( .A(n418), .B(n417), .Z(n450) );
  INV_X1 U478 ( .A(n450), .ZN(n419) );
  XOR2_X1 U479 ( .A(n420), .B(n419), .Z(n457) );
  NOR2_X1 U480 ( .A1(n522), .A2(n423), .ZN(n570) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n425) );
  XNOR2_X1 U482 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U484 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U485 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n437) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n467) );
  NAND2_X1 U494 ( .A1(n570), .A2(n467), .ZN(n440) );
  XOR2_X1 U495 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT65), .Z(n446) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(KEYINPUT86), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n452) );
  XOR2_X1 U502 ( .A(n450), .B(n449), .Z(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n538) );
  NAND2_X1 U504 ( .A1(n453), .A2(n538), .ZN(n566) );
  NOR2_X1 U505 ( .A1(n559), .A2(n566), .ZN(n456) );
  INV_X1 U506 ( .A(KEYINPUT58), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n538), .B(KEYINPUT87), .ZN(n460) );
  INV_X1 U508 ( .A(n457), .ZN(n524) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n524), .ZN(n465) );
  NAND2_X1 U510 ( .A1(n465), .A2(n522), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT98), .ZN(n532) );
  NOR2_X1 U512 ( .A1(n532), .A2(n536), .ZN(n459) );
  NAND2_X1 U513 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U514 ( .A(KEYINPUT99), .B(n461), .ZN(n475) );
  XNOR2_X1 U515 ( .A(KEYINPUT101), .B(KEYINPUT26), .ZN(n463) );
  NOR2_X1 U516 ( .A1(n538), .A2(n467), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U518 ( .A(KEYINPUT100), .B(n464), .Z(n569) );
  NAND2_X1 U519 ( .A1(n465), .A2(n569), .ZN(n470) );
  NAND2_X1 U520 ( .A1(n538), .A2(n524), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NAND2_X1 U523 ( .A1(n470), .A2(n469), .ZN(n472) );
  NAND2_X1 U524 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U525 ( .A(KEYINPUT102), .B(n473), .Z(n474) );
  NOR2_X1 U526 ( .A1(n475), .A2(n474), .ZN(n493) );
  NAND2_X1 U527 ( .A1(n559), .A2(n579), .ZN(n476) );
  XNOR2_X1 U528 ( .A(n476), .B(KEYINPUT16), .ZN(n477) );
  XNOR2_X1 U529 ( .A(n477), .B(KEYINPUT84), .ZN(n478) );
  NOR2_X1 U530 ( .A1(n493), .A2(n478), .ZN(n508) );
  NOR2_X1 U531 ( .A1(n571), .A2(n576), .ZN(n496) );
  NAND2_X1 U532 ( .A1(n508), .A2(n496), .ZN(n479) );
  XNOR2_X1 U533 ( .A(n479), .B(KEYINPUT103), .ZN(n490) );
  NAND2_X1 U534 ( .A1(n490), .A2(n522), .ZN(n483) );
  XOR2_X1 U535 ( .A(KEYINPUT34), .B(KEYINPUT106), .Z(n481) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(KEYINPUT105), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U539 ( .A(KEYINPUT104), .B(n484), .ZN(G1324GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n486) );
  NAND2_X1 U541 ( .A1(n490), .A2(n524), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U545 ( .A1(n490), .A2(n538), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT109), .Z(n492) );
  NAND2_X1 U548 ( .A1(n490), .A2(n536), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT110), .B(KEYINPUT39), .Z(n499) );
  NOR2_X1 U551 ( .A1(n585), .A2(n493), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n494), .A2(n567), .ZN(n495) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n495), .ZN(n521) );
  NAND2_X1 U554 ( .A1(n496), .A2(n521), .ZN(n497) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n497), .Z(n504) );
  NAND2_X1 U556 ( .A1(n522), .A2(n504), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n504), .A2(n524), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n538), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT111), .Z(n506) );
  NAND2_X1 U565 ( .A1(n536), .A2(n504), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  NOR2_X1 U567 ( .A1(n507), .A2(n562), .ZN(n520) );
  AND2_X1 U568 ( .A1(n508), .A2(n520), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n517), .A2(n522), .ZN(n512) );
  XOR2_X1 U570 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n510) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U574 ( .A(KEYINPUT112), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n517), .A2(n524), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT115), .Z(n516) );
  NAND2_X1 U578 ( .A1(n517), .A2(n538), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U581 ( .A1(n517), .A2(n536), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  AND2_X1 U583 ( .A1(n521), .A2(n520), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n529), .A2(n522), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n529), .A2(n524), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n527) );
  NAND2_X1 U589 ( .A1(n529), .A2(n538), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n536), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U596 ( .A(n534), .B(KEYINPUT119), .Z(n549) );
  INV_X1 U597 ( .A(n549), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n571), .A2(n545), .ZN(n539) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n562), .A2(n545), .ZN(n541) );
  XNOR2_X1 U603 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U606 ( .A1(n567), .A2(n545), .ZN(n543) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n559), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT121), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NAND2_X1 U613 ( .A1(n569), .A2(n549), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n571), .A2(n558), .ZN(n550) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n562), .A2(n558), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(KEYINPUT122), .B(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n567), .A2(n558), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT124), .B(n556), .Z(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n571), .A2(n566), .ZN(n561) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n566), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n584) );
  NOR2_X1 U636 ( .A1(n584), .A2(n571), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  INV_X1 U642 ( .A(n584), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n580), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

