//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G87), .B2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G68), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n220), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n211), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n210), .B(new_n214), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT12), .B1(new_n255), .B2(new_n221), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT74), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n253), .A2(KEYINPUT74), .A3(G13), .A4(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT12), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n260), .A2(new_n261), .A3(new_n225), .ZN(new_n262));
  INV_X1    g0062(.A(new_n260), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n207), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n221), .B1(new_n253), .B2(G20), .ZN(new_n267));
  AOI211_X1 g0067(.A(new_n256), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT73), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n208), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT73), .B1(G20), .B2(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n270), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n225), .A2(new_n208), .B1(new_n277), .B2(new_n215), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n265), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT11), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n280), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n268), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n289), .A2(KEYINPUT70), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT70), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(G1), .A2(G13), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G238), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G97), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G226), .A2(G1698), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n240), .B2(G1698), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT3), .B(G33), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n299), .B1(new_n305), .B2(new_n297), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n294), .A2(new_n306), .A3(KEYINPUT13), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n240), .A2(G1698), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G226), .B2(G1698), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n300), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n297), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n297), .A2(new_n298), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n315), .A2(new_n316), .B1(new_n317), .B2(G238), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n289), .A2(new_n291), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n289), .A2(KEYINPUT70), .A3(new_n291), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n308), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n307), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n283), .B1(G190), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n307), .B2(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT13), .B1(new_n294), .B2(new_n306), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n318), .A2(new_n323), .A3(new_n308), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT76), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT14), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(KEYINPUT76), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT77), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G169), .B1(new_n307), .B2(new_n324), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .A4(KEYINPUT14), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT78), .B(KEYINPUT14), .Z(new_n343));
  AOI22_X1  g0143(.A1(new_n325), .A2(G179), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n329), .B1(new_n345), .B2(new_n283), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT65), .B(G68), .ZN(new_n347));
  INV_X1    g0147(.A(G58), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n202), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n271), .A2(new_n272), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n349), .A2(G20), .B1(G159), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT79), .B1(new_n312), .B2(G33), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT79), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(new_n270), .A3(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n354), .A3(new_n313), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n356), .A3(new_n208), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n355), .B2(new_n208), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n351), .B(KEYINPUT16), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n201), .B1(new_n225), .B2(G58), .ZN(new_n362));
  INV_X1    g0162(.A(G159), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n362), .A2(new_n208), .B1(new_n363), .B2(new_n273), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n356), .A2(KEYINPUT80), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n304), .B2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n314), .A2(new_n208), .A3(new_n367), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n347), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n361), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n360), .A2(new_n372), .A3(new_n265), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT8), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G58), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n348), .A2(KEYINPUT8), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT71), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n265), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G1), .B2(new_n208), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n255), .B2(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n297), .A2(G232), .A3(new_n298), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n292), .B2(new_n293), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(G226), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(G1698), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n389), .A2(new_n352), .A3(new_n313), .A4(new_n354), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n297), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n330), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT81), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n388), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G223), .B2(G1698), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n391), .B1(new_n355), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n316), .ZN(new_n398));
  INV_X1    g0198(.A(G179), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n323), .A2(new_n398), .A3(new_n399), .A4(new_n385), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n393), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n394), .B1(new_n393), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n384), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT18), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n384), .B(new_n405), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(G200), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n386), .B2(new_n392), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n323), .A2(new_n398), .A3(new_n409), .A4(new_n385), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(new_n373), .A3(new_n383), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n411), .A2(new_n373), .A3(new_n383), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT17), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n404), .A2(new_n406), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n277), .B1(new_n376), .B2(new_n378), .ZN(new_n419));
  OAI21_X1  g0219(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n420));
  INV_X1    g0220(.A(G150), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n273), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n265), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  MUX2_X1   g0223(.A(new_n254), .B(new_n381), .S(G50), .Z(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G222), .A2(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G1698), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(G223), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n304), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n297), .B1(new_n314), .B2(new_n215), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n429), .A2(new_n430), .B1(new_n317), .B2(G226), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n323), .A3(new_n399), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n323), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n330), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n425), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n317), .A2(G244), .ZN(new_n436));
  NOR2_X1   g0236(.A1(G232), .A2(G1698), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n427), .A2(G238), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n304), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n316), .C1(G107), .C2(new_n304), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n323), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(new_n409), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(G200), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n266), .B(G77), .C1(G1), .C2(new_n208), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT15), .B(G87), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n375), .A2(new_n377), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n350), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n265), .B1(new_n215), .B2(new_n263), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n441), .A2(G179), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n444), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n441), .A2(new_n330), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT75), .B1(new_n433), .B2(new_n409), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(G200), .B2(new_n433), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n425), .A2(KEYINPUT9), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT9), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n423), .A2(new_n424), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT10), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT10), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n435), .B(new_n457), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n346), .A2(new_n418), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n208), .B1(new_n300), .B2(new_n471), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  INV_X1    g0275(.A(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(KEYINPUT84), .A3(new_n471), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n352), .A2(new_n354), .A3(new_n208), .A4(new_n313), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n478), .B(new_n479), .C1(new_n221), .C2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(new_n265), .B1(new_n445), .B2(new_n263), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G238), .A2(G1698), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n216), .B2(G1698), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(new_n352), .A3(new_n313), .A4(new_n354), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n297), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n284), .A2(new_n290), .A3(G1), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G250), .B1(new_n284), .B2(G1), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n316), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(G200), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n270), .B2(G1), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n253), .A2(KEYINPUT82), .A3(G33), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n496), .A2(new_n380), .A3(new_n254), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n216), .A2(G1698), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G238), .B2(G1698), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n486), .B1(new_n355), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n316), .ZN(new_n502));
  INV_X1    g0302(.A(new_n491), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(G190), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n482), .A2(new_n492), .A3(new_n498), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n472), .A2(new_n473), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n474), .A2(new_n477), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n479), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n480), .A2(new_n221), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n265), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n446), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n263), .A2(new_n445), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n330), .B1(new_n487), .B2(new_n491), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n502), .A2(new_n503), .A3(new_n399), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n215), .B1(new_n271), .B2(new_n272), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n520), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n519), .B1(new_n524), .B2(new_n208), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n217), .B1(new_n369), .B2(new_n370), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n265), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n496), .A2(new_n380), .A3(G97), .A4(new_n254), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n255), .A2(new_n521), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n216), .A2(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n352), .A2(new_n354), .A3(new_n313), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G250), .A2(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT4), .A2(G244), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G1698), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n304), .A2(new_n539), .B1(G33), .B2(G283), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n316), .ZN(new_n542));
  XNOR2_X1  g0342(.A(KEYINPUT5), .B(G41), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n284), .A2(G1), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n543), .A2(new_n544), .B1(new_n295), .B2(new_n296), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G257), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n543), .A2(new_n488), .A3(new_n297), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n542), .A2(new_n399), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n297), .B1(new_n536), .B2(new_n540), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n545), .A2(G257), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n550), .A2(new_n551), .A3(new_n547), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n532), .B(new_n549), .C1(G169), .C2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n542), .A2(G190), .A3(new_n546), .A4(new_n548), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT83), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n542), .A2(new_n546), .A3(new_n548), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G200), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n369), .A2(new_n370), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G107), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n521), .A2(new_n217), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n520), .B1(new_n560), .B2(new_n475), .ZN(new_n561));
  INV_X1    g0361(.A(new_n522), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n518), .B1(new_n563), .B2(G20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n530), .B1(new_n565), .B2(new_n265), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n541), .A2(new_n316), .B1(G257), .B2(new_n545), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(G190), .A4(new_n548), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n555), .A2(new_n557), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n517), .A2(new_n553), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n543), .A2(new_n544), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(G264), .A3(new_n297), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT85), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT85), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n545), .A2(new_n575), .A3(G264), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g0377(.A1(G250), .A2(G1698), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G257), .B2(new_n427), .ZN(new_n579));
  INV_X1    g0379(.A(G294), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n355), .A2(new_n579), .B1(new_n270), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n547), .B1(new_n581), .B2(new_n316), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(G179), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n547), .B1(G264), .B2(new_n545), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n316), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n330), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT22), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n208), .A2(G87), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n314), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n486), .A2(G20), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT23), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n208), .B2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n217), .A2(KEYINPUT23), .A3(G20), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n588), .A2(new_n476), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n480), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT24), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n352), .A2(new_n354), .A3(new_n313), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n208), .A3(new_n597), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n590), .A4(new_n595), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n380), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n497), .A2(G107), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n254), .A2(G107), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT25), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n584), .A2(new_n587), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(new_n604), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n265), .ZN(new_n612));
  INV_X1    g0412(.A(new_n609), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n585), .A2(new_n409), .A3(new_n586), .ZN(new_n614));
  AOI21_X1  g0414(.A(G200), .B1(new_n577), .B2(new_n582), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n218), .A2(G1698), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G257), .B2(G1698), .ZN(new_n619));
  INV_X1    g0419(.A(G303), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n355), .A2(new_n619), .B1(new_n620), .B2(new_n304), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n316), .ZN(new_n622));
  OR2_X1    g0422(.A1(KEYINPUT5), .A2(G41), .ZN(new_n623));
  NAND2_X1  g0423(.A1(KEYINPUT5), .A2(G41), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n295), .B2(new_n296), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n545), .A2(G270), .B1(new_n488), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G200), .ZN(new_n628));
  INV_X1    g0428(.A(G116), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n263), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n260), .A2(G116), .A3(new_n380), .A4(new_n496), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n264), .A2(new_n207), .B1(G20), .B2(new_n629), .ZN(new_n632));
  AOI21_X1  g0432(.A(G20), .B1(G33), .B2(G283), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G33), .B2(new_n521), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT20), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n632), .A2(new_n634), .A3(KEYINPUT20), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n630), .B(new_n631), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n628), .B(new_n638), .C1(new_n409), .C2(new_n627), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n622), .A2(new_n626), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(G179), .A3(new_n637), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n330), .B1(new_n622), .B2(new_n626), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n642), .A2(new_n643), .A3(new_n637), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n642), .B2(new_n637), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n639), .B(new_n641), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n617), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n469), .A2(new_n571), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT86), .Z(G372));
  AND2_X1   g0449(.A1(new_n404), .A2(new_n406), .ZN(new_n650));
  INV_X1    g0450(.A(new_n456), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n345), .A2(new_n283), .B1(new_n328), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n416), .A2(new_n414), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n465), .A2(new_n467), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n435), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n469), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n658));
  INV_X1    g0458(.A(new_n587), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n612), .A2(new_n613), .B1(new_n659), .B2(new_n583), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n616), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n517), .A2(new_n570), .A3(new_n553), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n516), .ZN(new_n664));
  AOI21_X1  g0464(.A(G169), .B1(new_n567), .B2(new_n548), .ZN(new_n665));
  NOR4_X1   g0465(.A1(new_n550), .A2(new_n551), .A3(G179), .A4(new_n547), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n566), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n517), .A2(new_n667), .A3(KEYINPUT26), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n505), .A2(new_n516), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n553), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n664), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n656), .B1(new_n657), .B2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n253), .A2(new_n208), .A3(G13), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT27), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n253), .A3(new_n208), .A4(G13), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(G213), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  XOR2_X1   g0481(.A(KEYINPUT88), .B(G343), .Z(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n638), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n658), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n646), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n685), .B1(new_n612), .B2(new_n613), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n691), .A2(new_n617), .B1(new_n610), .B2(new_n685), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n658), .A2(new_n685), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(new_n617), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n660), .A2(new_n685), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n696), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n477), .A2(G116), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n212), .A2(new_n288), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n205), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(new_n685), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n663), .B2(new_n672), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI211_X1 g0511(.A(KEYINPUT29), .B(new_n708), .C1(new_n663), .C2(new_n672), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n487), .A2(new_n491), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n640), .A2(new_n567), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n716), .B2(new_n583), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n502), .A2(new_n503), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n627), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n584), .A2(new_n719), .A3(KEYINPUT30), .A4(new_n567), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n627), .A2(new_n718), .A3(new_n399), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n567), .A2(new_n548), .B1(new_n577), .B2(new_n582), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n577), .A2(new_n582), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n556), .A2(new_n724), .A3(KEYINPUT91), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n717), .B(new_n720), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n708), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n647), .A2(new_n571), .A3(new_n685), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n713), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n707), .B1(new_n735), .B2(G1), .ZN(G364));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n253), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n704), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n690), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n688), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n304), .A2(new_n212), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n212), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n355), .A2(new_n212), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n285), .A2(new_n287), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n205), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n251), .B2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n747), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n295), .B1(new_n208), .B2(G169), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT93), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT93), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n742), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n208), .A2(new_n399), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n409), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n208), .B1(new_n768), .B2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n766), .A2(new_n767), .B1(new_n770), .B2(G294), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G326), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n208), .A2(new_n409), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n407), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n304), .B1(new_n778), .B2(G303), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n771), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n208), .A2(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n768), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n783), .A2(G283), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n399), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT94), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n781), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n781), .B2(new_n788), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n780), .B(new_n790), .C1(G311), .C2(new_n795), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n304), .B1(new_n782), .B2(new_n217), .C1(new_n476), .C2(new_n777), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n769), .A2(new_n521), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G68), .B2(new_n766), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT97), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n785), .A2(G159), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n798), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n772), .A2(new_n274), .B1(new_n789), .B2(new_n348), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n795), .B2(G77), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT95), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n796), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT98), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n757), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n763), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n760), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n688), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n744), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n811), .A2(new_n759), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n742), .B1(new_n818), .B2(G77), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT99), .ZN(new_n820));
  INV_X1    g0620(.A(new_n789), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G294), .A2(new_n821), .B1(new_n783), .B2(G87), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n823), .B2(new_n784), .C1(new_n629), .C2(new_n794), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n314), .B1(new_n777), .B2(new_n217), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n799), .B1(G283), .B2(new_n766), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n620), .B2(new_n772), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n773), .A2(G137), .B1(new_n821), .B2(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n831), .B1(new_n421), .B2(new_n765), .C1(new_n363), .C2(new_n794), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT102), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n777), .A2(new_n274), .B1(new_n782), .B2(new_n221), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n601), .B1(new_n348), .B2(new_n769), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G132), .C2(new_n785), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n830), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n820), .B1(new_n840), .B2(new_n811), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(KEYINPUT103), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n842), .A2(KEYINPUT103), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT104), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n456), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n453), .A2(KEYINPUT104), .A3(new_n454), .A4(new_n455), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n846), .A2(new_n452), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n708), .A2(new_n454), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n848), .A2(new_n849), .B1(new_n651), .B2(new_n708), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n843), .B(new_n844), .C1(new_n758), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT26), .B1(new_n517), .B2(new_n667), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n670), .A2(new_n553), .A3(new_n669), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n516), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n661), .A2(new_n662), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n685), .B(new_n848), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n849), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n708), .A2(new_n651), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n709), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n860), .A2(new_n733), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n742), .B1(new_n860), .B2(new_n733), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n851), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n738), .A2(new_n253), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n345), .A2(new_n283), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n708), .A2(new_n283), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n328), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n283), .B(new_n708), .C1(new_n345), .C2(new_n329), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n846), .A2(new_n847), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n685), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n856), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n681), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n373), .B2(new_n383), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n415), .A2(new_n876), .A3(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n403), .A2(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT105), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n384), .B(new_n879), .C1(new_n401), .C2(new_n402), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n360), .A2(new_n265), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT7), .B1(new_n601), .B2(G20), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(G68), .A3(new_n357), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT16), .B1(new_n884), .B2(new_n351), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n383), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n401), .B2(new_n402), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n412), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n886), .A2(new_n681), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n881), .A2(new_n890), .B1(new_n417), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n881), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n417), .A2(new_n889), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n871), .B(new_n874), .C1(new_n892), .C2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n650), .B2(new_n681), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT108), .ZN(new_n898));
  XNOR2_X1  g0698(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n881), .A2(KEYINPUT107), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT107), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n877), .A2(new_n878), .A3(new_n901), .A4(new_n880), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n415), .A2(new_n876), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n403), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n900), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n417), .A2(new_n876), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n898), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT39), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n881), .A2(KEYINPUT107), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(new_n902), .B1(new_n417), .B2(new_n876), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n913), .B(KEYINPUT108), .C1(new_n915), .C2(new_n899), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n892), .B2(new_n895), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n867), .A2(new_n708), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n897), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n469), .B1(new_n711), .B2(new_n712), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n656), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n920), .B(new_n922), .Z(new_n923));
  INV_X1    g0723(.A(G330), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT31), .B1(new_n726), .B2(new_n708), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n850), .B1(new_n927), .B2(new_n730), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n871), .A2(new_n928), .A3(KEYINPUT40), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n909), .B1(new_n915), .B2(new_n899), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT109), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n906), .A2(new_n907), .ZN(new_n933));
  INV_X1    g0733(.A(new_n899), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n895), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n871), .A2(new_n928), .A3(KEYINPUT40), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n871), .B(new_n928), .C1(new_n892), .C2(new_n895), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n931), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n469), .A2(new_n732), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n924), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n866), .B1(new_n923), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n923), .B2(new_n943), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n563), .A2(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n563), .A2(KEYINPUT35), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(G116), .A3(new_n209), .A4(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n206), .B(G77), .C1(new_n348), .C2(new_n347), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(G50), .B2(new_n221), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(G1), .A3(new_n737), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n945), .A2(new_n949), .A3(new_n952), .ZN(G367));
  OAI211_X1 g0753(.A(new_n570), .B(new_n553), .C1(new_n685), .C2(new_n566), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n708), .A2(new_n667), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(new_n695), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n954), .A2(new_n610), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n708), .B1(new_n960), .B2(new_n553), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n958), .B2(KEYINPUT42), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n685), .B1(new_n482), .B2(new_n498), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n517), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n959), .A2(new_n962), .B1(KEYINPUT43), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n693), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n956), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n704), .B(KEYINPUT41), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n701), .A2(new_n956), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT45), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n701), .A2(new_n956), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n969), .ZN(new_n978));
  INV_X1    g0778(.A(new_n694), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n695), .B1(new_n692), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n689), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n734), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n974), .A2(new_n976), .A3(new_n693), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n978), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n972), .B1(new_n986), .B2(new_n735), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n971), .B1(new_n987), .B2(new_n740), .ZN(new_n988));
  INV_X1    g0788(.A(new_n749), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n238), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n761), .B1(new_n212), .B2(new_n445), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n742), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n795), .A2(G50), .ZN(new_n993));
  INV_X1    g0793(.A(G137), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n782), .A2(new_n215), .B1(new_n784), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G58), .B2(new_n778), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n304), .B1(new_n789), .B2(new_n421), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G159), .B2(new_n766), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n773), .A2(G143), .B1(new_n770), .B2(G68), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n993), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n782), .A2(new_n521), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G303), .B2(new_n821), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n1003), .B2(new_n784), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT46), .B1(new_n777), .B2(new_n629), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n629), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G283), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n794), .A2(new_n1008), .B1(new_n217), .B2(new_n769), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT111), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n355), .B1(new_n765), .B2(new_n580), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G311), .B2(new_n773), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1009), .A2(KEYINPUT111), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1000), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT47), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n811), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n992), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n965), .B2(new_n814), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n988), .A2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n734), .A2(new_n981), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n982), .A2(new_n741), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n981), .A2(new_n739), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n692), .A2(new_n814), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n745), .A2(new_n703), .B1(G107), .B2(new_n212), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT112), .Z(new_n1028));
  INV_X1    g0828(.A(new_n243), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n750), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n448), .A2(new_n274), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n703), .B(new_n284), .C1(new_n221), .C2(new_n215), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n989), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1028), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n742), .B1(new_n1036), .B2(new_n762), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n789), .A2(new_n274), .B1(new_n784), .B2(new_n421), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1001), .B(new_n1038), .C1(G77), .C2(new_n778), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n769), .A2(new_n445), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n355), .B(new_n1040), .C1(G159), .C2(new_n773), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n379), .A2(new_n766), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n795), .A2(G68), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n783), .A2(G116), .B1(new_n785), .B2(G326), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n777), .A2(new_n580), .B1(new_n769), .B2(new_n1008), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n766), .A2(G311), .B1(new_n821), .B2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n787), .B2(new_n772), .C1(new_n620), .C2(new_n794), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n355), .B(new_n1045), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1044), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1037), .B1(new_n1055), .B2(new_n757), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1025), .B1(new_n1026), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1024), .A2(new_n1057), .ZN(G393));
  NAND2_X1  g0858(.A1(new_n978), .A2(new_n984), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n982), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n741), .A3(new_n986), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n978), .A2(new_n740), .A3(new_n984), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT113), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n777), .A2(new_n1008), .B1(new_n784), .B2(new_n787), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n304), .B(new_n1064), .C1(G107), .C2(new_n783), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n772), .A2(new_n1003), .B1(new_n789), .B2(new_n823), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n795), .A2(G294), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n766), .A2(G303), .B1(new_n770), .B2(G116), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n772), .A2(new_n421), .B1(new_n789), .B2(new_n363), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n769), .A2(new_n215), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n355), .B(new_n1073), .C1(G50), .C2(new_n766), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n795), .A2(new_n448), .ZN(new_n1075));
  INV_X1    g0875(.A(G143), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n782), .A2(new_n476), .B1(new_n784), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n225), .B2(new_n778), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n811), .B1(new_n1070), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n989), .A2(new_n247), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n761), .B1(new_n521), .B2(new_n212), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n742), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n956), .B2(new_n814), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1062), .A2(new_n1063), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1063), .B1(new_n1062), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1061), .B1(new_n1086), .B2(new_n1087), .ZN(G390));
  NAND3_X1  g0888(.A1(new_n469), .A2(G330), .A3(new_n732), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n921), .A2(new_n656), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n871), .A2(new_n928), .A3(G330), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n732), .A2(G330), .A3(new_n859), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n869), .A3(new_n870), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n874), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n871), .A2(new_n874), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n919), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n912), .A2(new_n916), .A3(new_n1100), .A4(new_n917), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n930), .A2(new_n1099), .A3(new_n1098), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n1091), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1091), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1105));
  OAI211_X1 g0905(.A(KEYINPUT114), .B(new_n1097), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1091), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1097), .A2(KEYINPUT114), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1103), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1106), .A2(new_n741), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n740), .A3(new_n1103), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n742), .B1(new_n818), .B2(new_n379), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n777), .A2(new_n421), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT53), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1115), .A2(new_n1116), .B1(new_n1117), .B2(new_n772), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1116), .B2(new_n1115), .ZN(new_n1119));
  INV_X1    g0919(.A(G132), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n789), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n304), .B1(new_n782), .B2(new_n274), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G125), .C2(new_n785), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n794), .A2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n766), .A2(G137), .B1(new_n770), .B2(G159), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1119), .A2(new_n1123), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n304), .B(new_n1073), .C1(G87), .C2(new_n778), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n795), .A2(G97), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G107), .A2(new_n766), .B1(new_n773), .B2(G283), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n782), .A2(new_n221), .B1(new_n784), .B2(new_n580), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G116), .B2(new_n821), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1114), .B1(new_n1134), .B2(new_n757), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n918), .B2(new_n759), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1112), .A2(new_n1113), .A3(new_n1136), .ZN(G378));
  OAI21_X1  g0937(.A(new_n742), .B1(new_n818), .B2(G50), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n355), .A2(new_n288), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1139), .B(new_n274), .C1(G33), .C2(G41), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n794), .A2(new_n445), .B1(new_n521), .B2(new_n765), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT115), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G107), .A2(new_n821), .B1(new_n785), .B2(G283), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n348), .B2(new_n782), .C1(new_n215), .C2(new_n777), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n772), .A2(new_n629), .B1(new_n769), .B2(new_n221), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n1142), .A2(new_n1139), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1140), .B1(new_n1146), .B2(KEYINPUT58), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT116), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n794), .A2(new_n994), .B1(new_n1120), .B2(new_n765), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT117), .Z(new_n1150));
  AOI22_X1  g0950(.A1(new_n773), .A2(G125), .B1(new_n770), .B2(G150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n777), .A2(new_n1124), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G128), .B2(new_n821), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n363), .B2(new_n782), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1156), .B2(KEYINPUT59), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1157), .A2(new_n1160), .B1(KEYINPUT58), .B2(new_n1146), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1148), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1138), .B1(new_n1162), .B2(new_n757), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n435), .B1(new_n465), .B2(new_n467), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n425), .A2(new_n681), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1164), .B(new_n1165), .Z(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1163), .B1(new_n1168), .B2(new_n759), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT120), .Z(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n920), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n931), .A2(new_n937), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n924), .B1(new_n939), .B2(new_n938), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n1168), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1168), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n935), .A2(new_n936), .A3(new_n932), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT109), .B1(new_n929), .B2(new_n930), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1168), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1173), .A2(new_n1174), .A3(new_n1168), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n920), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1171), .B1(new_n1185), .B2(new_n740), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1109), .A2(new_n1103), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1090), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1175), .A2(new_n1176), .A3(new_n1172), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n920), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(KEYINPUT57), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n741), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1186), .B1(new_n1194), .B2(new_n1195), .ZN(G375));
  OAI21_X1  g0996(.A(new_n742), .B1(new_n818), .B2(G68), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n304), .B(new_n1040), .C1(G77), .C2(new_n783), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n795), .A2(G107), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G116), .A2(new_n766), .B1(new_n773), .B2(G294), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n777), .A2(new_n521), .B1(new_n784), .B2(new_n620), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G283), .B2(new_n821), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n794), .A2(new_n421), .B1(new_n274), .B2(new_n769), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT122), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n601), .B1(new_n772), .B2(new_n1120), .C1(new_n765), .C2(new_n1124), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n777), .A2(new_n363), .B1(new_n782), .B2(new_n348), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n789), .A2(new_n994), .B1(new_n784), .B2(new_n1117), .ZN(new_n1208));
  OR3_X1    g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1197), .B1(new_n1210), .B2(new_n757), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n871), .B2(new_n759), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1187), .B2(new_n739), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n874), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n921), .A2(new_n656), .A3(new_n1089), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n972), .B(KEYINPUT121), .Z(new_n1220));
  NAND3_X1  g1020(.A1(new_n1097), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1214), .A2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT123), .Z(G381));
  NAND3_X1  g1023(.A1(new_n1024), .A2(new_n816), .A3(new_n1057), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1224), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G378), .A2(new_n1225), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n682), .A2(G213), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT124), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(G213), .A3(new_n1231), .ZN(G409));
  NAND2_X1  g1032(.A1(new_n1230), .A2(G2897), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1217), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1219), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1187), .A2(KEYINPUT60), .A3(new_n1217), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n741), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT125), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n704), .B1(new_n1241), .B2(new_n1219), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT125), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1238), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1245), .B2(new_n1214), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n864), .B(new_n1213), .C1(new_n1240), .C2(new_n1244), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1234), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1243), .B1(new_n1242), .B2(new_n1238), .ZN(new_n1249));
  AND4_X1   g1049(.A1(new_n1243), .A2(new_n1237), .A3(new_n741), .A4(new_n1238), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1214), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n864), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1245), .A2(G384), .A3(new_n1214), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1233), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G378), .B(new_n1186), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1185), .A2(new_n740), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1170), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1185), .A2(new_n1190), .A3(new_n1220), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1228), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1230), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G387), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G390), .A2(new_n988), .A3(new_n1021), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n816), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(KEYINPUT126), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT126), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1273), .A2(new_n1269), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1264), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1230), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1277), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1265), .A2(new_n1275), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1280), .A2(new_n1283), .A3(new_n1277), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1280), .B2(new_n1255), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1283), .B1(new_n1280), .B2(new_n1277), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1284), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT127), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1273), .A2(new_n1269), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1270), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1282), .B1(new_n1288), .B2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1228), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1257), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1277), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1278), .A2(new_n1297), .A3(new_n1257), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1275), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G402));
endmodule


