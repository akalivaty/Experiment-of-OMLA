//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT70), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G127gat), .B2(new_n202), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n203), .A2(new_n205), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n203), .A2(KEYINPUT70), .ZN(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n224), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n230), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT69), .B1(new_n230), .B2(new_n231), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(G190gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT28), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT27), .B1(new_n234), .B2(KEYINPUT68), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n242), .C1(KEYINPUT68), .C2(new_n237), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n232), .A2(new_n233), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n227), .A3(new_n228), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n224), .A3(KEYINPUT25), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(G183gat), .A3(G190gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G183gat), .B(G190gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n251), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n234), .A2(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n238), .A2(G183gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n252), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT66), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n261), .B(new_n252), .C1(new_n253), .C2(new_n251), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n248), .A2(new_n247), .B1(new_n221), .B2(new_n223), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n255), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n219), .B1(new_n245), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT72), .B(new_n219), .C1(new_n245), .C2(new_n266), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n221), .A2(new_n223), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n229), .A2(new_n225), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n231), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n230), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n276));
  INV_X1    g075(.A(new_n244), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n219), .ZN(new_n279));
  INV_X1    g078(.A(new_n265), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n249), .A2(new_n224), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(KEYINPUT66), .B2(new_n254), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n282), .B2(new_n262), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n278), .B(new_n279), .C1(new_n283), .C2(new_n255), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT71), .ZN(new_n285));
  INV_X1    g084(.A(new_n266), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n279), .A4(new_n278), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n269), .A2(new_n270), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G227gat), .A2(G233gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n290), .B(KEYINPUT64), .Z(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT34), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n291), .A2(KEYINPUT34), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  XOR2_X1   g094(.A(G15gat), .B(G43gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT73), .ZN(new_n297));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n300), .B2(new_n299), .ZN(new_n302));
  INV_X1    g101(.A(new_n292), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT32), .B(new_n302), .C1(new_n289), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n269), .A2(new_n270), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n288), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT33), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n294), .B(new_n304), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n306), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n292), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT32), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n295), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n316), .A3(new_n299), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n294), .A4(new_n304), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n304), .B1(new_n310), .B2(new_n308), .ZN(new_n320));
  INV_X1    g119(.A(new_n294), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n312), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT36), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n322), .A2(KEYINPUT36), .A3(new_n311), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G1gat), .B(G29gat), .Z(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  OR2_X1    g132(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n335));
  INV_X1    g134(.A(G141gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G148gat), .ZN(new_n337));
  INV_X1    g136(.A(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(G141gat), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n334), .B(new_n335), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT78), .B1(new_n336), .B2(G148gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(new_n338), .A3(G141gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n336), .A2(G148gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n341), .B1(new_n350), .B2(KEYINPUT2), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n340), .A2(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n353));
  NAND3_X1  g152(.A1(new_n279), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n351), .ZN(new_n355));
  XNOR2_X1  g154(.A(G141gat), .B(G148gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n344), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n214), .A2(new_n218), .A3(new_n355), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n355), .A2(new_n358), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n214), .A2(KEYINPUT79), .A3(new_n218), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT79), .B1(new_n214), .B2(new_n218), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n366), .B(new_n368), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n359), .A2(new_n353), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n352), .A2(new_n360), .A3(new_n214), .A4(new_n218), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n375), .A3(new_n364), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n364), .B1(new_n377), .B2(new_n359), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(KEYINPUT5), .C1(new_n378), .C2(KEYINPUT81), .ZN(new_n379));
  INV_X1    g178(.A(new_n359), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n219), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n214), .A2(KEYINPUT79), .A3(new_n218), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n380), .B1(new_n384), .B2(new_n367), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n385), .A2(new_n386), .A3(new_n364), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n333), .B(new_n372), .C1(new_n379), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n385), .B2(new_n364), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n378), .A2(KEYINPUT81), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT5), .A4(new_n376), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n333), .B1(new_n393), .B2(new_n372), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT91), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(KEYINPUT6), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n372), .B1(new_n379), .B2(new_n387), .ZN(new_n397));
  INV_X1    g196(.A(new_n333), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n389), .A4(new_n388), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT38), .ZN(new_n403));
  AND2_X1   g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n245), .B2(new_n266), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n278), .B(new_n405), .C1(new_n283), .C2(new_n255), .ZN(new_n409));
  XNOR2_X1  g208(.A(G197gat), .B(G204gat), .ZN(new_n410));
  INV_X1    g209(.A(G211gat), .ZN(new_n411));
  INV_X1    g210(.A(G218gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(KEYINPUT22), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G211gat), .B(G218gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n408), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n408), .B2(new_n409), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT37), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT37), .B1(new_n418), .B2(new_n419), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT76), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n427), .B2(KEYINPUT93), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT93), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n429), .A3(new_n426), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n403), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n409), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n416), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n408), .A2(new_n409), .A3(new_n417), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n425), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(new_n403), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n420), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n419), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n418), .A2(KEYINPUT92), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n435), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n402), .A2(new_n431), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT85), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT31), .B(G50gat), .Z(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(KEYINPUT86), .B2(G22gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(G22gat), .B2(new_n448), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n417), .B1(new_n366), .B2(new_n406), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n365), .B1(new_n416), .B2(KEYINPUT29), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n367), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n450), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G228gat), .A2(G233gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n455), .B(KEYINPUT87), .Z(new_n456));
  XNOR2_X1  g255(.A(new_n454), .B(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n434), .A4(new_n425), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n426), .B1(new_n418), .B2(new_n419), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n459), .A2(KEYINPUT88), .A3(new_n460), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n371), .A2(new_n354), .A3(new_n361), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  INV_X1    g267(.A(new_n364), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n333), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n377), .A2(new_n364), .A3(new_n359), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT39), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n473), .A2(new_n474), .B1(new_n467), .B2(new_n469), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(KEYINPUT89), .A3(KEYINPUT39), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n477), .A2(KEYINPUT40), .B1(new_n398), .B2(new_n397), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n467), .A2(new_n469), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n364), .B1(new_n362), .B2(new_n371), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n398), .B1(new_n483), .B2(new_n468), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI211_X1 g286(.A(KEYINPUT90), .B(KEYINPUT40), .C1(new_n482), .C2(new_n484), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n478), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n457), .B1(new_n466), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n444), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n399), .A2(new_n389), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n397), .B2(new_n398), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(new_n390), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n394), .A2(new_n495), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n499), .B2(new_n462), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n389), .B(new_n388), .C1(new_n394), .C2(new_n495), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n399), .A2(KEYINPUT83), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n396), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n462), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT84), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n457), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n328), .A2(new_n492), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n322), .A2(new_n311), .A3(new_n457), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n500), .A3(new_n505), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT94), .B(KEYINPUT35), .Z(new_n513));
  NAND4_X1  g312(.A1(new_n402), .A2(new_n466), .A3(new_n457), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n323), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT98), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT9), .ZN(new_n521));
  NAND2_X1  g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n520), .B2(new_n519), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(KEYINPUT96), .A2(G71gat), .A3(G78gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT100), .B(G64gat), .Z(new_n534));
  NAND2_X1  g333(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n522), .B1(new_n527), .B2(new_n521), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT101), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G127gat), .B(G155gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT20), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G183gat), .B(G211gat), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(G1gat), .B2(new_n551), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(G8gat), .Z(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n539), .B2(new_n540), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT102), .B(KEYINPUT19), .Z(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n556), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n550), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n548), .A2(new_n560), .A3(new_n549), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT15), .ZN(new_n565));
  OR2_X1    g364(.A1(G43gat), .A2(G50gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G43gat), .A2(G50gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT95), .B(G43gat), .Z(new_n569));
  OAI211_X1 g368(.A(new_n565), .B(new_n567), .C1(new_n569), .C2(G50gat), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT14), .B(G29gat), .Z(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(G36gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n568), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n568), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT17), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT105), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n579), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n591), .A2(KEYINPUT106), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(KEYINPUT106), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n577), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT41), .ZN(new_n598));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT103), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n595), .B(new_n597), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n598), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT104), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n602), .ZN(new_n608));
  AND4_X1   g407(.A1(KEYINPUT107), .A2(new_n603), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(KEYINPUT107), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n603), .B2(new_n608), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n564), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n578), .A2(new_n555), .ZN(new_n615));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n555), .A2(new_n575), .A3(new_n576), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT18), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n555), .B(new_n577), .Z(new_n620));
  XOR2_X1   g419(.A(new_n616), .B(KEYINPUT13), .Z(new_n621));
  AOI22_X1  g420(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n615), .A2(new_n617), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(KEYINPUT18), .A3(new_n616), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT11), .B(G169gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n622), .B2(new_n624), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n594), .A2(new_n539), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n591), .B(KEYINPUT106), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n533), .A2(new_n538), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT108), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n588), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n588), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n589), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n635), .A2(new_n642), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G120gat), .B(G148gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT109), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n648), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n634), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n614), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n518), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n499), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g465(.A1(new_n663), .A2(new_n466), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G8gat), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT111), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT42), .B1(new_n667), .B2(KEYINPUT110), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(G1325gat));
  AOI21_X1  g476(.A(new_n326), .B1(new_n323), .B2(new_n324), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT112), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n663), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n323), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n663), .B2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n663), .A2(new_n457), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NOR2_X1   g485(.A1(new_n564), .A2(new_n661), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n518), .A2(new_n612), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n571), .A3(new_n499), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n457), .B1(new_n500), .B2(new_n505), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n491), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n693), .A2(new_n328), .B1(new_n512), .B2(new_n516), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n694), .B2(new_n613), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n518), .A2(KEYINPUT44), .A3(new_n612), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n687), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n503), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n690), .A2(new_n699), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n698), .B2(new_n466), .ZN(new_n701));
  INV_X1    g500(.A(G36gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n466), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n705), .A3(new_n706), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n697), .A2(new_n678), .A3(new_n687), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n569), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n323), .A2(new_n569), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n688), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n678), .B(KEYINPUT112), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n713), .A3(new_n687), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n714), .A2(new_n569), .B1(new_n688), .B2(new_n710), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n715), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g515(.A1(new_n695), .A2(new_n696), .A3(new_n507), .A4(new_n687), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n688), .A2(new_n719), .A3(new_n507), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT48), .B1(new_n721), .B2(KEYINPUT113), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  AOI211_X1 g523(.A(new_n723), .B(new_n724), .C1(new_n718), .C2(new_n720), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n725), .ZN(G1331gat));
  NOR3_X1   g525(.A1(new_n614), .A2(new_n660), .A3(new_n634), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT114), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n518), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n499), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n518), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n466), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n323), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n729), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G71gat), .B1(new_n732), .B2(new_n680), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n732), .A2(new_n457), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT115), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  NOR3_X1   g546(.A1(new_n564), .A2(new_n660), .A3(new_n634), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n697), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n503), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n564), .A2(new_n634), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n678), .A2(new_n692), .A3(new_n491), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n515), .B1(KEYINPUT35), .B2(new_n511), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n612), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n518), .A2(KEYINPUT51), .A3(new_n612), .A4(new_n751), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n660), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n584), .A3(new_n499), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT116), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n750), .B1(new_n759), .B2(new_n762), .ZN(G1336gat));
  NAND4_X1  g562(.A1(new_n695), .A2(new_n696), .A3(new_n703), .A4(new_n748), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n660), .A2(new_n466), .A3(G92gat), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT117), .B1(new_n758), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768));
  INV_X1    g567(.A(new_n766), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n768), .B(new_n769), .C1(new_n756), .C2(new_n757), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n765), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(new_n758), .B2(new_n766), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n764), .A2(G92gat), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n771), .A2(new_n772), .B1(new_n776), .B2(new_n777), .ZN(G1337gat));
  OR4_X1    g577(.A1(G99gat), .A2(new_n759), .A3(new_n323), .A4(new_n660), .ZN(new_n779));
  OAI21_X1  g578(.A(G99gat), .B1(new_n749), .B2(new_n680), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(G1338gat));
  NOR2_X1   g580(.A1(new_n457), .A2(G106gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n758), .A2(new_n760), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n695), .A2(new_n696), .A3(new_n507), .A4(new_n748), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT119), .B(G106gat), .Z(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g587(.A(new_n564), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n644), .A2(new_n650), .A3(new_n645), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n648), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n650), .B1(new_n644), .B2(new_n645), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n658), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n659), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(new_n791), .B2(new_n794), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT120), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n791), .A2(new_n794), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n659), .A4(new_n795), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n634), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n623), .A2(new_n616), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n620), .A2(new_n621), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n628), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n630), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n660), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n612), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n609), .A2(new_n808), .A3(new_n611), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n798), .A3(new_n803), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n789), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n564), .A2(new_n613), .A3(new_n660), .A4(new_n633), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n703), .A2(new_n503), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n739), .A3(new_n457), .A4(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n209), .A3(new_n633), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n510), .A3(new_n634), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(new_n209), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n819), .B2(new_n660), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n510), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n760), .A2(new_n207), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT121), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n825), .B2(new_n827), .ZN(G1341gat));
  OAI21_X1  g627(.A(G127gat), .B1(new_n819), .B2(new_n789), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n564), .A2(new_n204), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n825), .B2(new_n830), .ZN(G1342gat));
  NAND2_X1  g630(.A1(new_n612), .A2(new_n202), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n825), .A2(KEYINPUT56), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n819), .B2(new_n613), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT56), .B1(new_n825), .B2(new_n832), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  INV_X1    g635(.A(new_n816), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n801), .A2(new_n659), .A3(new_n795), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n633), .B1(new_n838), .B2(KEYINPUT122), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n796), .A2(KEYINPUT122), .A3(new_n797), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n809), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n813), .B1(new_n841), .B2(new_n612), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n837), .B1(new_n842), .B2(new_n789), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT57), .B1(new_n843), .B2(new_n457), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n457), .B1(new_n815), .B2(new_n816), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n678), .A2(new_n503), .A3(new_n703), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n844), .A2(new_n847), .A3(new_n634), .A4(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(G141gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n680), .A2(new_n507), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT123), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(KEYINPUT123), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n821), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n633), .A2(G141gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT58), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n849), .A2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n859), .B(new_n860), .C1(new_n854), .C2(new_n856), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(G1344gat));
  INV_X1    g661(.A(new_n854), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n338), .A3(new_n760), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT59), .B(new_n338), .C1(new_n865), .C2(new_n760), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n845), .A2(new_n846), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n841), .A2(new_n612), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n613), .A2(new_n808), .A3(new_n838), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n789), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n816), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n457), .A2(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n868), .A2(new_n760), .A3(new_n874), .A4(new_n848), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n864), .B1(new_n866), .B2(new_n876), .ZN(G1345gat));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n844), .A2(new_n847), .A3(new_n564), .A4(new_n848), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(G155gat), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n789), .A2(G155gat), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n854), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(G155gat), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(KEYINPUT124), .C1(new_n854), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1346gat));
  AOI21_X1  g686(.A(G162gat), .B1(new_n863), .B2(new_n612), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n612), .A2(G162gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n865), .B2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n499), .A2(new_n466), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n815), .B2(new_n816), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n510), .ZN(new_n894));
  AOI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n634), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n323), .A2(new_n507), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n227), .A3(new_n633), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n898), .ZN(G1348gat));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n228), .A3(new_n760), .ZN(new_n900));
  OAI21_X1  g699(.A(G176gat), .B1(new_n897), .B2(new_n660), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1349gat));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n897), .B2(new_n789), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n893), .A2(KEYINPUT125), .A3(new_n564), .A4(new_n896), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(G183gat), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n564), .A2(new_n235), .A3(new_n237), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n894), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT60), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n906), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n894), .A2(new_n238), .A3(new_n612), .ZN(new_n915));
  OAI21_X1  g714(.A(G190gat), .B1(new_n897), .B2(new_n613), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(KEYINPUT61), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(KEYINPUT61), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n713), .A2(new_n892), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n868), .A2(new_n874), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(G197gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(new_n633), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n920), .A2(new_n845), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n634), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n923), .B1(new_n928), .B2(new_n922), .ZN(G1352gat));
  INV_X1    g728(.A(G204gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n924), .A2(new_n930), .A3(new_n760), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT62), .ZN(new_n932));
  OAI21_X1  g731(.A(G204gat), .B1(new_n921), .B2(new_n660), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G1353gat));
  NAND4_X1  g734(.A1(new_n868), .A2(new_n564), .A3(new_n874), .A4(new_n920), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n926), .A2(new_n927), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n564), .A2(new_n411), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n938), .A2(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n921), .B2(new_n613), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n612), .A2(new_n412), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n940), .B2(new_n944), .ZN(G1355gat));
endmodule


