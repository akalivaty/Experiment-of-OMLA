//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340;
  OR2_X1    g0000(.A1(KEYINPUT64), .A2(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(KEYINPUT64), .A2(G50), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n202), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n207), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n217), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  INV_X1    g0041(.A(KEYINPUT3), .ZN(new_n242));
  INV_X1    g0042(.A(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n246), .A2(G222), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n246), .A2(G223), .A3(G1698), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n248), .B(new_n249), .C1(new_n250), .C2(new_n246), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(G274), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n259), .B(KEYINPUT66), .C1(new_n260), .C2(new_n263), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n253), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G179), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(new_n214), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n261), .A2(G20), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G50), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n215), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n204), .A2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n204), .A2(new_n288), .A3(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n275), .A2(new_n214), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n274), .B(new_n279), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n253), .A2(new_n266), .A3(new_n267), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n270), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  AOI22_X1  g0098(.A1(G190), .A2(new_n268), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n293), .A2(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n294), .A2(new_n303), .A3(G200), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n294), .B2(G200), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n279), .A2(new_n274), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n287), .A2(new_n289), .ZN(new_n310));
  INV_X1    g0110(.A(new_n285), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n309), .B1(new_n312), .B2(new_n291), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n313), .A2(KEYINPUT9), .B1(new_n294), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n300), .ZN(new_n316));
  INV_X1    g0116(.A(new_n305), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n294), .A2(new_n303), .A3(G200), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n308), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n297), .B1(new_n307), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G58), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n202), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n283), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n244), .A2(new_n215), .A3(new_n245), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n244), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n245), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n332), .A2(KEYINPUT71), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT71), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(new_n331), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n329), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n328), .B1(new_n339), .B2(new_n327), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n291), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(new_n292), .A3(new_n271), .A4(new_n278), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n280), .A2(new_n272), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n322), .A2(KEYINPUT8), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n322), .A2(KEYINPUT8), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n278), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n346), .B(new_n343), .C1(new_n350), .C2(new_n276), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n258), .A2(G232), .A3(new_n262), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n259), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n260), .A2(G1698), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n357), .B1(G223), .B2(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n314), .B(new_n356), .C1(new_n362), .C2(new_n258), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n258), .B1(new_n360), .B2(new_n361), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n355), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n341), .A2(new_n342), .A3(new_n353), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT74), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n347), .A2(new_n352), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n332), .A2(KEYINPUT71), .A3(new_n333), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(G68), .A3(new_n336), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n292), .B1(new_n372), .B2(new_n329), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n373), .B2(new_n340), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n342), .A4(new_n367), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n341), .A2(new_n353), .A3(new_n367), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT73), .B1(new_n378), .B2(KEYINPUT17), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n378), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n365), .A2(new_n355), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n295), .B2(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT18), .B1(new_n385), .B2(new_n374), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n341), .A2(new_n353), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n384), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n263), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G244), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n259), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT68), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n246), .A2(G232), .A3(new_n247), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n246), .A2(G238), .A3(G1698), .ZN(new_n399));
  INV_X1    g0199(.A(G107), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n398), .B(new_n399), .C1(new_n400), .C2(new_n246), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n252), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(KEYINPUT68), .A3(new_n259), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n269), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n344), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT15), .B(G87), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n281), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n291), .B1(new_n250), .B2(new_n272), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n278), .A2(G77), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n276), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT69), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n295), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(G200), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n413), .B(new_n409), .C1(new_n415), .C2(new_n314), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n272), .A2(new_n323), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT12), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n323), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n250), .B2(new_n281), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n277), .A2(G68), .A3(new_n278), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT11), .B1(new_n427), .B2(new_n291), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n246), .A2(G232), .A3(G1698), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n246), .A2(G226), .A3(new_n247), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G97), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n252), .ZN(new_n438));
  INV_X1    g0238(.A(G274), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n252), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(G238), .A2(new_n393), .B1(new_n440), .B2(new_n256), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT13), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n438), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(G179), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n445), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n438), .B2(new_n441), .ZN(new_n448));
  OAI21_X1  g0248(.A(G169), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n449), .B2(KEYINPUT14), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(new_n445), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G169), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n433), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G200), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n443), .A2(G190), .A3(new_n445), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n432), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n423), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n321), .A2(new_n392), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT75), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n243), .B2(G1), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n261), .A2(KEYINPUT75), .A3(G33), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n277), .A2(new_n463), .A3(G116), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n272), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n275), .A2(new_n214), .B1(G20), .B2(new_n465), .ZN(new_n468));
  AOI21_X1  g0268(.A(G20), .B1(G33), .B2(G283), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n243), .A2(G97), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT81), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT81), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT20), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n261), .B(G45), .C1(new_n254), .C2(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT77), .B1(new_n480), .B2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT77), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n254), .A3(KEYINPUT5), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT78), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT78), .B1(new_n481), .B2(new_n483), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n479), .B(new_n440), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G264), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n487));
  OAI211_X1 g0287(.A(G257), .B(new_n247), .C1(new_n358), .C2(new_n359), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n244), .A2(G303), .A3(new_n245), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n252), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n481), .A2(new_n483), .ZN(new_n492));
  OAI211_X1 g0292(.A(G270), .B(new_n258), .C1(new_n492), .C2(new_n478), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n486), .A2(new_n491), .A3(G179), .A4(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n477), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n486), .A2(new_n491), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G169), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n498), .B2(new_n477), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n499), .B2(KEYINPUT21), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n358), .A2(new_n359), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n215), .A3(G87), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n508));
  INV_X1    g0308(.A(G87), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(KEYINPUT83), .A3(G20), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n246), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G20), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT23), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n215), .B2(G107), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n400), .A2(KEYINPUT23), .A3(G20), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n507), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n291), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G13), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G1), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G20), .A3(new_n400), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(KEYINPUT85), .A3(KEYINPUT25), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT85), .B(KEYINPUT25), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n277), .A2(new_n463), .A3(KEYINPUT76), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n461), .A2(new_n462), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n276), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(G107), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G257), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n535));
  OAI211_X1 g0335(.A(G250), .B(new_n247), .C1(new_n358), .C2(new_n359), .ZN(new_n536));
  INV_X1    g0336(.A(G294), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n243), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n252), .ZN(new_n539));
  OAI211_X1 g0339(.A(G264), .B(new_n258), .C1(new_n492), .C2(new_n478), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n486), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G169), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT86), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(new_n486), .A3(G179), .A4(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n544), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n534), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n496), .B(new_n549), .C1(new_n498), .C2(new_n477), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n500), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n541), .A2(new_n314), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n541), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n521), .A3(new_n533), .A4(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G244), .B(new_n247), .C1(new_n358), .C2(new_n359), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n246), .A2(KEYINPUT4), .A3(G244), .A4(new_n247), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G283), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n246), .A2(G250), .A3(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n252), .ZN(new_n562));
  INV_X1    g0362(.A(new_n492), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n252), .B1(new_n563), .B2(new_n479), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G257), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n486), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n295), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  AND2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n400), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n573), .A2(new_n215), .B1(new_n250), .B2(new_n284), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n400), .B1(new_n332), .B2(new_n333), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n291), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n272), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n528), .A2(G97), .A3(new_n531), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n561), .A2(new_n252), .B1(new_n564), .B2(G257), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n269), .A3(new_n486), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n567), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n566), .A2(G200), .ZN(new_n584));
  INV_X1    g0384(.A(new_n575), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n571), .A2(new_n572), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(G20), .B1(G77), .B2(new_n283), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n292), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(new_n578), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n581), .A2(G190), .A3(new_n486), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n584), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n554), .A2(new_n583), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n497), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n477), .B1(new_n595), .B2(new_n364), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n497), .A2(new_n314), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n407), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n528), .A2(new_n531), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n215), .B1(new_n436), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n570), .A2(new_n509), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n215), .B(G68), .C1(new_n358), .C2(new_n359), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n281), .B2(new_n577), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n291), .B1(new_n272), .B2(new_n407), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  INV_X1    g0411(.A(G250), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n255), .B2(G1), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n261), .A2(new_n439), .A3(G45), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n258), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(G244), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n617));
  OAI211_X1 g0417(.A(G238), .B(new_n247), .C1(new_n358), .C2(new_n359), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n512), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n252), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(new_n295), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n269), .B(new_n616), .C1(new_n619), .C2(new_n252), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n611), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(G179), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(KEYINPUT79), .C1(new_n295), .C2(new_n620), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n610), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(G190), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT80), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n528), .A2(G87), .A3(new_n531), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n608), .C1(new_n620), .C2(new_n364), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT80), .B1(new_n620), .B2(G190), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n598), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n551), .A2(new_n594), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n459), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT87), .ZN(G372));
  NAND3_X1  g0437(.A1(new_n500), .A2(new_n548), .A3(new_n550), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n630), .A2(new_n608), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n619), .A2(new_n252), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n615), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n627), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n609), .B1(new_n621), .B2(new_n622), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(KEYINPUT88), .A3(new_n644), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n594), .A2(new_n638), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n644), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n567), .A2(new_n582), .A3(new_n580), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n643), .A2(KEYINPUT88), .A3(new_n644), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT88), .B1(new_n643), .B2(new_n644), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n626), .A2(new_n583), .A3(new_n633), .ZN(new_n657));
  XOR2_X1   g0457(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n652), .A2(new_n656), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n459), .ZN(new_n662));
  INV_X1    g0462(.A(new_n297), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n452), .A2(new_n451), .A3(G169), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n446), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n666), .A2(new_n433), .B1(new_n418), .B2(new_n457), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n378), .A2(KEYINPUT17), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT73), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n378), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(new_n369), .B2(new_n376), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n391), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n307), .A2(new_n320), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n663), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n662), .A2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n500), .A2(new_n550), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n523), .A2(new_n215), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n523), .A2(new_n680), .A3(new_n215), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(G213), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n477), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n677), .B(new_n685), .Z(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n598), .ZN(new_n687));
  INV_X1    g0487(.A(new_n684), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n548), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n534), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n554), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n548), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n687), .A2(G330), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n677), .A2(new_n684), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n208), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n603), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n212), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(new_n684), .C1(new_n651), .C2(new_n660), .ZN(new_n709));
  INV_X1    g0509(.A(new_n644), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n654), .A2(new_n655), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n593), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n712), .B2(new_n638), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n656), .A2(new_n652), .B1(new_n657), .B2(new_n659), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n688), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n709), .B1(new_n715), .B2(new_n708), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n566), .A2(new_n717), .A3(new_n541), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n566), .B2(new_n541), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n497), .A2(new_n269), .A3(new_n641), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n497), .A2(new_n641), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n546), .A3(new_n581), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n546), .A3(KEYINPUT30), .A4(new_n581), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n688), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n635), .A2(new_n684), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n688), .C1(new_n721), .C2(new_n727), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT92), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n716), .B1(G330), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n707), .B1(new_n737), .B2(G1), .ZN(G364));
  NAND2_X1  g0538(.A1(new_n687), .A2(G330), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n522), .A2(G20), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT93), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n261), .A3(new_n702), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n687), .A2(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n686), .B2(new_n598), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n246), .A2(new_n208), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n208), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n237), .A2(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n701), .A2(new_n246), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n255), .B2(new_n213), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n214), .B1(G20), .B2(new_n295), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n751), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n744), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(G20), .A2(G179), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(new_n314), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n323), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n215), .A2(G179), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT32), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n765), .A2(new_n314), .A3(new_n364), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n273), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G87), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n774), .B2(new_n773), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n766), .A2(new_n770), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n364), .A2(G190), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n765), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n246), .B1(new_n250), .B2(new_n783), .C1(new_n786), .C2(new_n322), .ZN(new_n787));
  OR4_X1    g0587(.A1(new_n768), .A2(new_n778), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(G20), .B1(new_n784), .B2(G179), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT95), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G97), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n769), .A2(new_n314), .A3(G200), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT94), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT94), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n400), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n767), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G303), .A2(new_n780), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n783), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n246), .B1(new_n804), .B2(G311), .ZN(new_n805));
  INV_X1    g0605(.A(new_n771), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G329), .B1(new_n785), .B2(G322), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n776), .A2(G326), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n803), .A2(new_n805), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n537), .A2(new_n793), .B1(new_n799), .B2(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n788), .A2(new_n800), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n764), .B1(new_n812), .B2(new_n761), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n748), .B1(new_n752), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n661), .A2(new_n684), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n418), .A2(new_n684), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n688), .A2(new_n414), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n420), .B2(new_n421), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n417), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n821), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n823), .B(new_n684), .C1(new_n651), .C2(new_n660), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n736), .A2(G330), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n744), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n761), .A2(new_n749), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT96), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n744), .B1(new_n830), .B2(G77), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n780), .A2(G107), .B1(G303), .B2(new_n776), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n810), .B2(new_n767), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n504), .B1(new_n786), .B2(new_n537), .ZN(new_n834));
  INV_X1    g0634(.A(G311), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n771), .A2(new_n835), .B1(new_n783), .B2(new_n465), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n799), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G87), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n795), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n246), .B1(new_n771), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n799), .A2(new_n323), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n843), .C1(G50), .C2(new_n780), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n322), .B2(new_n793), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n804), .A2(G159), .B1(G143), .B2(new_n785), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n777), .C1(new_n282), .C2(new_n767), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT34), .Z(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n831), .B1(new_n850), .B2(new_n761), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n823), .B2(new_n750), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n828), .A2(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n586), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n586), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n216), .A4(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OR3_X1    g0658(.A1(new_n212), .A2(new_n250), .A3(new_n324), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n201), .A2(new_n203), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(G68), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n261), .B(G13), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n338), .A2(new_n291), .ZN(new_n865));
  INV_X1    g0665(.A(new_n327), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT16), .B1(new_n372), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n346), .B(new_n345), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(new_n683), .B1(new_n374), .B2(new_n367), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n384), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n378), .B1(new_n385), .B2(new_n374), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n387), .A2(new_n683), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT99), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n387), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n871), .B1(new_n864), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n868), .A2(new_n683), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT98), .B1(new_n392), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT98), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n883), .B(new_n880), .C1(new_n381), .C2(new_n391), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n879), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT38), .B(new_n879), .C1(new_n882), .C2(new_n884), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n670), .A2(new_n671), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n390), .B1(new_n891), .B2(new_n377), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n883), .B1(new_n892), .B2(new_n880), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT98), .B(new_n881), .C1(new_n672), .C2(new_n390), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n886), .B(new_n878), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n877), .A2(new_n864), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n877), .A2(new_n864), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n875), .A2(new_n876), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n392), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n890), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n666), .A2(new_n433), .A3(new_n684), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n889), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n391), .A2(new_n683), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n887), .A2(new_n888), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n433), .A2(new_n688), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n454), .A2(new_n457), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n457), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n433), .B(new_n688), .C1(new_n666), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n824), .B2(new_n817), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n906), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT100), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n905), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n905), .B2(new_n915), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n321), .A2(new_n458), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n892), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n583), .B1(new_n647), .B2(new_n648), .ZN(new_n922));
  INV_X1    g0722(.A(new_n633), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n623), .A2(new_n625), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n653), .B(new_n923), .C1(new_n610), .C2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n922), .A2(KEYINPUT26), .B1(new_n925), .B2(new_n658), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n684), .B1(new_n651), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT29), .ZN(new_n928));
  AOI211_X1 g0728(.A(KEYINPUT101), .B(new_n921), .C1(new_n928), .C2(new_n709), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT101), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n716), .B2(new_n459), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n675), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n919), .B(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(G330), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n551), .A2(new_n594), .A3(new_n634), .A4(new_n684), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n730), .A3(new_n733), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n821), .B1(new_n909), .B2(new_n911), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n893), .A2(new_n894), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n940), .B2(new_n879), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n941), .B2(new_n895), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT40), .ZN(new_n943));
  INV_X1    g0743(.A(new_n900), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n896), .A2(new_n897), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n886), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n888), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT102), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT40), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT102), .B1(new_n936), .B2(new_n937), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n942), .A2(new_n943), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n459), .A2(new_n936), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n934), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n933), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n261), .B2(new_n740), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n933), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n863), .B1(new_n958), .B2(new_n959), .ZN(G367));
  OAI211_X1 g0760(.A(new_n583), .B(new_n592), .C1(new_n590), .C2(new_n684), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n653), .A2(new_n688), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n698), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n684), .A2(new_n639), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n649), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n644), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n583), .B1(new_n961), .B2(new_n548), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n684), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n966), .A2(new_n973), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n970), .B(KEYINPUT43), .Z(new_n976));
  AOI22_X1  g0776(.A1(new_n974), .A2(KEYINPUT103), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n974), .A2(KEYINPUT103), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n695), .A2(new_n964), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(new_n977), .B2(new_n978), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n702), .B(new_n983), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n699), .A2(new_n963), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT106), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n699), .A2(new_n963), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n699), .A2(new_n963), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n699), .B2(new_n963), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n695), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n697), .B(new_n693), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n739), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n737), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n992), .A2(new_n695), .A3(new_n996), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n985), .B1(new_n1004), .B2(new_n737), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n743), .A2(new_n261), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n982), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n838), .A2(G97), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1010), .B(new_n504), .C1(new_n1011), .C2(new_n771), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT107), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n804), .A2(G283), .B1(G303), .B2(new_n785), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n537), .B2(new_n767), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G311), .B2(new_n776), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n780), .A2(G116), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT46), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n400), .C2(new_n793), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n1014), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n793), .A2(new_n323), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G150), .B2(new_n785), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT108), .Z(new_n1025));
  OAI221_X1 g0825(.A(new_n246), .B1(new_n771), .B2(new_n847), .C1(new_n860), .C2(new_n783), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n780), .A2(G58), .B1(G143), .B2(new_n776), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n772), .B2(new_n767), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(G77), .C2(new_n838), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1022), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT109), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n761), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n968), .A2(new_n751), .A3(new_n969), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n233), .A2(new_n757), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n763), .B1(new_n701), .B2(new_n599), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n745), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n1009), .A2(KEYINPUT110), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT110), .B1(new_n1009), .B2(new_n1039), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n693), .A2(new_n751), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n753), .A2(new_n704), .B1(G107), .B2(new_n208), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n758), .B1(new_n230), .B2(G45), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n255), .B1(new_n323), .B2(new_n250), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n704), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT111), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT50), .B1(new_n344), .B2(new_n273), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n344), .A2(KEYINPUT50), .A3(new_n273), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1045), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1044), .B(new_n744), .C1(new_n763), .C2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT112), .B(G150), .Z(new_n1056));
  OAI22_X1  g0856(.A1(new_n786), .A2(new_n273), .B1(new_n1056), .B2(new_n771), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n504), .B(new_n1057), .C1(G68), .C2(new_n804), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n780), .A2(G77), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n280), .B2(new_n767), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G159), .B2(new_n776), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n794), .A2(new_n599), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1061), .A3(new_n1010), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n804), .A2(G303), .B1(G317), .B2(new_n785), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n776), .A2(G322), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n835), .C2(new_n767), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT113), .Z(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT48), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT48), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n794), .A2(G283), .B1(G294), .B2(new_n780), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n838), .A2(G116), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n246), .B1(new_n806), .B2(G326), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1063), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1055), .B1(new_n1079), .B2(new_n761), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1001), .A2(new_n702), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1000), .A2(new_n737), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(G393));
  INV_X1    g0884(.A(new_n1003), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1085), .A2(new_n997), .A3(new_n1006), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n964), .A2(new_n751), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n762), .B1(new_n577), .B2(new_n208), .C1(new_n240), .C2(new_n758), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n744), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n786), .A2(new_n835), .B1(new_n777), .B2(new_n1011), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT52), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n794), .A2(G116), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n504), .B1(new_n783), .B2(new_n537), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G322), .B2(new_n806), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G283), .A2(new_n780), .B1(new_n801), .B2(G303), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n799), .C2(new_n400), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n860), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1098), .A2(new_n801), .B1(new_n780), .B2(G68), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n806), .A2(G143), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n504), .B1(new_n804), .B2(new_n344), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n839), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n794), .A2(G77), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n785), .A2(G159), .B1(new_n776), .B2(G150), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT51), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(KEYINPUT51), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1093), .A2(new_n1097), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1089), .B1(new_n1108), .B2(new_n761), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1086), .B1(new_n1087), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1001), .B1(new_n1085), .B2(new_n997), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n1004), .A3(new_n702), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(G390));
  INV_X1    g0913(.A(new_n820), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n817), .B1(new_n927), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n912), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n947), .A3(new_n903), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n821), .A2(new_n934), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n732), .B2(new_n735), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n912), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT39), .B1(new_n888), .B2(new_n946), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n941), .A2(new_n895), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(KEYINPUT39), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n914), .A2(new_n904), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1117), .B(new_n1121), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n936), .A2(new_n912), .A3(new_n1118), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n889), .B2(new_n902), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1117), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1126), .A2(new_n1131), .A3(new_n1007), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n744), .B1(new_n830), .B2(new_n344), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1056), .A2(new_n779), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT53), .Z(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n246), .B1(new_n783), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n786), .A2(new_n841), .B1(new_n771), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n777), .A2(new_n1140), .B1(new_n847), .B2(new_n767), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n772), .B2(new_n793), .C1(new_n860), .C2(new_n799), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1103), .B1(new_n465), .B2(new_n786), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT117), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n781), .B1(new_n400), .B2(new_n767), .C1(new_n810), .C2(new_n777), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n504), .B1(new_n783), .B2(new_n577), .C1(new_n537), .C2(new_n771), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n843), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1133), .B1(new_n1149), .B2(new_n761), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1124), .B2(new_n750), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1132), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n459), .A2(G330), .A3(new_n936), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT114), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT114), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n459), .A2(new_n1156), .A3(G330), .A4(new_n936), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n675), .B(new_n1158), .C1(new_n929), .C2(new_n931), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1127), .B1(new_n1120), .B2(new_n912), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n824), .A2(new_n817), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n912), .B1(new_n936), .B2(new_n1118), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1115), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1160), .A2(new_n1161), .B1(new_n1163), .B2(new_n1121), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n889), .A2(new_n902), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1125), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1127), .B1(new_n1168), .B2(new_n1117), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1121), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1129), .A2(new_n1130), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT115), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(KEYINPUT115), .A3(new_n1165), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1126), .A2(new_n1131), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n702), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT116), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT116), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1183), .B(new_n1180), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1153), .B1(new_n1182), .B2(new_n1184), .ZN(G378));
  NAND3_X1  g0985(.A1(new_n905), .A2(new_n915), .A3(new_n916), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n905), .A2(new_n915), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT100), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n951), .A2(new_n947), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n938), .B1(new_n887), .B2(new_n888), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(G330), .C1(new_n1190), .C2(KEYINPUT40), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n293), .A2(new_n683), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n321), .B(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1195));
  XOR2_X1   g0995(.A(new_n1194), .B(new_n1195), .Z(new_n1196));
  NOR2_X1   g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1196), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n952), .B2(G330), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1186), .B(new_n1188), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT123), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n952), .A2(G330), .A3(new_n1198), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n917), .C2(new_n918), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1159), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1179), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n919), .B(KEYINPUT123), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1210), .B1(new_n1179), .B2(new_n1206), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n703), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1205), .A2(new_n1007), .A3(new_n1208), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1196), .A2(new_n749), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n829), .A2(new_n860), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n838), .A2(G58), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT119), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G41), .B(new_n246), .C1(new_n804), .C2(new_n599), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n400), .B2(new_n786), .C1(new_n810), .C2(new_n771), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1059), .B1(new_n577), .B2(new_n767), .C1(new_n465), .C2(new_n777), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1220), .A2(new_n1023), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n777), .A2(new_n1138), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n786), .A2(new_n1140), .B1(new_n783), .B2(new_n847), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(G132), .C2(new_n801), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n779), .A2(new_n1136), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT120), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n282), .C2(new_n793), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n243), .A2(new_n254), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT118), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G124), .B2(new_n806), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n799), .B2(new_n772), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT121), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1232), .A2(new_n1233), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1235), .B(new_n273), .C1(G41), .C2(new_n246), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1225), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n745), .B(new_n1218), .C1(new_n1242), .C2(new_n761), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1217), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1216), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1215), .A2(new_n1246), .ZN(G375));
  NOR2_X1   g1047(.A1(new_n1164), .A2(new_n1006), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n913), .A2(new_n749), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n744), .B1(new_n830), .B2(G68), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n786), .A2(new_n810), .B1(new_n783), .B2(new_n400), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n246), .B(new_n1251), .C1(G303), .C2(new_n806), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n838), .A2(G77), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n779), .A2(new_n577), .B1(new_n767), .B2(new_n465), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G294), .B2(new_n776), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1062), .A4(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n786), .A2(new_n847), .B1(new_n771), .B2(new_n1140), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n504), .B(new_n1257), .C1(G150), .C2(new_n804), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n794), .A2(G50), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n776), .A2(G132), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1136), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G159), .A2(new_n780), .B1(new_n801), .B2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .A4(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1256), .B1(new_n1220), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1250), .B1(new_n1264), .B2(new_n761), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1248), .B1(new_n1249), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1165), .A2(new_n984), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(G381));
  OR4_X1    g1069(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(G387), .A2(G381), .A3(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G375), .B(KEYINPUT124), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1173), .B(new_n1178), .C1(new_n1126), .C2(new_n1131), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT115), .B1(new_n1175), .B2(new_n1165), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1181), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1153), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1271), .A2(new_n1272), .A3(new_n1277), .ZN(G407));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(G343), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(new_n1281), .A3(G213), .ZN(G409));
  NAND3_X1  g1082(.A1(G378), .A2(new_n1215), .A3(new_n1246), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1205), .A2(new_n984), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1212), .A2(new_n1007), .B1(new_n1217), .B2(new_n1243), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1276), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1280), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1268), .B1(new_n1165), .B2(KEYINPUT60), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n1164), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n702), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1266), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G384), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1266), .C1(new_n1289), .C2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1294), .A2(KEYINPUT125), .A3(new_n1295), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1288), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G393), .B(new_n814), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1008), .A2(G390), .A3(new_n1038), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n1008), .B2(new_n1038), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1305), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT127), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1311), .B(new_n1305), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1307), .A2(new_n1305), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1042), .B2(G390), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT61), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1280), .A2(G2897), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1298), .A2(new_n1299), .A3(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1296), .A2(G2897), .A3(new_n1280), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(KEYINPUT126), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1319), .A2(new_n1323), .A3(new_n1320), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1245), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1286), .B1(new_n1325), .B2(G378), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1322), .B(new_n1324), .C1(new_n1280), .C2(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1304), .A2(new_n1316), .A3(new_n1317), .A4(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1288), .B2(new_n1321), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1288), .B2(new_n1301), .ZN(new_n1332));
  NOR4_X1   g1132(.A1(new_n1326), .A2(KEYINPUT62), .A3(new_n1280), .A4(new_n1300), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1330), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1328), .B1(new_n1334), .B2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1277), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1300), .B1(new_n1337), .B2(new_n1283), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1337), .A2(new_n1283), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1296), .B2(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1335), .ZN(G402));
endmodule


