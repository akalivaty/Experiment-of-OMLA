//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT93), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n204), .A3(G1gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT94), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n212), .A2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(new_n223), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n216), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n233), .A3(new_n214), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n211), .A2(new_n233), .A3(new_n214), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n211), .B2(new_n214), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n229), .A2(new_n230), .A3(new_n223), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(new_n227), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n228), .A2(KEYINPUT17), .A3(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n235), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n202), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n228), .B(new_n231), .C1(new_n236), .C2(new_n237), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n235), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n245), .B(KEYINPUT13), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n217), .A2(new_n234), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n242), .A3(new_n241), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n245), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G169gat), .B(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n247), .A2(new_n252), .A3(new_n255), .A4(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(KEYINPUT95), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(G227gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n281), .A2(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT64), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n286), .A2(G169gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n287), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n282), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n284), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n286), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n296), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n309), .A2(KEYINPUT25), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n278), .A2(new_n302), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n292), .ZN(new_n316));
  OR3_X1    g115(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT68), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n303), .A2(new_n317), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n292), .B1(new_n312), .B2(new_n313), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT28), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n316), .A2(new_n322), .A3(new_n288), .A4(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329));
  INV_X1    g128(.A(G113gat), .ZN(new_n330));
  INV_X1    g129(.A(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT69), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G120gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n331), .A2(G113gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n328), .B(new_n329), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338));
  INV_X1    g137(.A(new_n329), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(KEYINPUT1), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n337), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n337), .B2(new_n341), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n311), .A2(new_n327), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n302), .A2(new_n278), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n307), .A2(new_n310), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n337), .A2(new_n338), .A3(new_n341), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .A4(new_n326), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n277), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n273), .B1(new_n352), .B2(KEYINPUT33), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n344), .A2(new_n351), .ZN(new_n357));
  AOI221_X4 g156(.A(new_n354), .B1(KEYINPUT33), .B2(new_n273), .C1(new_n357), .C2(new_n276), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n344), .A2(new_n351), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n344), .B2(new_n351), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n362), .A2(new_n363), .A3(new_n276), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n365));
  OAI21_X1  g164(.A(KEYINPUT74), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n344), .A2(new_n351), .A3(new_n361), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n277), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n370));
  INV_X1    g169(.A(new_n365), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n357), .A2(KEYINPUT34), .A3(new_n276), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n360), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g175(.A(KEYINPUT75), .B(new_n374), .C1(new_n366), .C2(new_n372), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n359), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT76), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  INV_X1    g181(.A(G211gat), .ZN(new_n383));
  INV_X1    g182(.A(G218gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n379), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT77), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n379), .A2(new_n381), .A3(new_n390), .A4(new_n385), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G226gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n275), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n311), .B2(new_n327), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n347), .B2(new_n326), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n393), .B(new_n396), .C1(new_n397), .C2(new_n395), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT79), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n393), .B(KEYINPUT78), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n397), .A2(new_n395), .ZN(new_n401));
  INV_X1    g200(.A(new_n396), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n395), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n311), .A2(new_n327), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(KEYINPUT29), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n393), .A4(new_n396), .ZN(new_n408));
  XOR2_X1   g207(.A(G8gat), .B(G36gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G64gat), .ZN(new_n410));
  INV_X1    g209(.A(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n399), .A2(new_n403), .A3(new_n408), .A4(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n414), .A2(KEYINPUT30), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(KEYINPUT30), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n403), .A3(new_n408), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n417), .A2(KEYINPUT80), .A3(new_n412), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT80), .B1(new_n417), .B2(new_n412), .ZN(new_n419));
  OAI22_X1  g218(.A1(new_n415), .A2(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424));
  OR2_X1    g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(KEYINPUT2), .ZN(new_n426));
  XOR2_X1   g225(.A(G141gat), .B(G148gat), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT81), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n424), .A3(new_n425), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n432), .A2(new_n435), .A3(new_n341), .A4(new_n337), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n423), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n431), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT81), .B1(new_n426), .B2(new_n427), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT3), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n432), .A2(new_n443), .A3(new_n435), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n348), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n441), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(new_n349), .A3(KEYINPUT4), .A4(new_n350), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n348), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n436), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n423), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT0), .B(G57gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(G85gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  OR2_X1    g256(.A1(new_n436), .A2(new_n437), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n349), .A2(new_n350), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n437), .B1(new_n459), .B2(new_n441), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n452), .A2(new_n423), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n445), .A4(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n453), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n457), .B1(new_n453), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n421), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n421), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n420), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n375), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n373), .A2(new_n360), .A3(new_n375), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n356), .B2(new_n358), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n357), .A2(new_n276), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT32), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n479), .A3(new_n273), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n353), .A2(new_n355), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT71), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n472), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G22gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(G228gat), .A2(G233gat), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n386), .A2(new_n380), .B1(new_n389), .B2(new_n391), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT85), .B1(new_n487), .B2(KEYINPUT29), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n393), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n491), .A3(new_n443), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n441), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n444), .A2(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n400), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n486), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n486), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n393), .B1(new_n444), .B2(new_n490), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n389), .A2(new_n391), .B1(new_n388), .B2(new_n386), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n490), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT84), .B1(new_n499), .B2(KEYINPUT29), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n443), .ZN(new_n504));
  AOI211_X1 g303(.A(new_n497), .B(new_n498), .C1(new_n504), .C2(new_n441), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n485), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT86), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n441), .ZN(new_n508));
  INV_X1    g307(.A(new_n498), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n486), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n492), .A2(new_n441), .B1(new_n400), .B2(new_n494), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n510), .B(G22gat), .C1(new_n511), .C2(new_n486), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G78gat), .B(G106gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT31), .ZN(new_n515));
  INV_X1    g314(.A(G50gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n507), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n506), .B(new_n512), .C1(KEYINPUT86), .C2(new_n517), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n378), .A2(new_n468), .A3(new_n484), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n376), .A2(new_n377), .A3(new_n359), .ZN(new_n528));
  INV_X1    g327(.A(new_n359), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n472), .B2(new_n473), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n472), .A2(new_n473), .A3(new_n529), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n378), .A2(KEYINPUT89), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(new_n521), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n468), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n525), .B(new_n526), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n484), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT36), .B1(new_n538), .B2(new_n530), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n378), .A2(new_n540), .A3(new_n532), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n521), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n458), .A2(new_n460), .A3(new_n445), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n423), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n547), .B(KEYINPUT39), .C1(new_n423), .C2(new_n450), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT39), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n549), .A3(new_n423), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n457), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT40), .ZN(new_n552));
  INV_X1    g351(.A(new_n464), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n420), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT87), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n406), .A2(new_n396), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n556), .A2(KEYINPUT88), .A3(new_n400), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n400), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT88), .B1(new_n556), .B2(new_n487), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n557), .B(KEYINPUT37), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n417), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT38), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n412), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n417), .B(KEYINPUT37), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT38), .B1(new_n565), .B2(new_n413), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n564), .A2(new_n566), .A3(new_n467), .A4(new_n414), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n420), .A3(new_n568), .A4(new_n553), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n555), .A2(new_n567), .A3(new_n521), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n543), .A2(new_n545), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n270), .B1(new_n537), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(G71gat), .ZN(new_n575));
  INV_X1    g374(.A(G78gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT9), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT96), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(KEYINPUT9), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584));
  AOI21_X1  g383(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n253), .A2(new_n383), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n383), .B1(new_n253), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n586), .A3(new_n589), .ZN(new_n594));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT20), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n592), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n592), .B2(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT19), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT97), .B(G183gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n598), .B2(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  OR2_X1    g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT99), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(G99gat), .A3(G106gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n617), .A3(KEYINPUT8), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n610), .B(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n620), .A2(new_n232), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n619), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n610), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n242), .A3(new_n241), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n625), .A3(new_n292), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n292), .B1(new_n622), .B2(new_n625), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n627), .A2(new_n628), .A3(new_n384), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(G190gat), .ZN(new_n631));
  AOI21_X1  g430(.A(G218gat), .B1(new_n631), .B2(new_n626), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n608), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT98), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n384), .B1(new_n627), .B2(new_n628), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n631), .A2(G218gat), .A3(new_n626), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT101), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n608), .B(new_n637), .C1(new_n629), .C2(new_n632), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n607), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n585), .A2(new_n610), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n610), .B1(new_n585), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n623), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n585), .A2(new_n610), .ZN(new_n650));
  AOI211_X1 g449(.A(KEYINPUT102), .B(new_n578), .C1(new_n583), .C2(new_n584), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n650), .B(new_n619), .C1(new_n651), .C2(new_n610), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT10), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n620), .A2(KEYINPUT10), .A3(new_n585), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G230gat), .ZN(new_n656));
  OAI22_X1  g455(.A1(new_n653), .A2(new_n655), .B1(new_n656), .B2(new_n275), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n275), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n649), .A2(new_n658), .A3(new_n652), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n284), .ZN(new_n662));
  INV_X1    g461(.A(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n657), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n572), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n467), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(new_n206), .ZN(G1324gat));
  INV_X1    g472(.A(new_n420), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n208), .A2(new_n213), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n680), .B(new_n681), .C1(new_n213), .C2(new_n675), .ZN(G1325gat));
  INV_X1    g481(.A(new_n670), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n531), .A2(new_n533), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n543), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(G15gat), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n670), .A2(new_n521), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n607), .A2(new_n644), .A3(new_n668), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI211_X1 g494(.A(new_n270), .B(new_n695), .C1(new_n537), .C2(new_n571), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n671), .A2(G29gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n537), .A2(new_n571), .ZN(new_n699));
  INV_X1    g498(.A(new_n270), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n697), .A4(new_n694), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(KEYINPUT103), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n692), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n693), .A3(new_n697), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(KEYINPUT103), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT104), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT104), .B1(new_n605), .B2(new_n606), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n266), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n712), .A3(new_n668), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n644), .A2(KEYINPUT44), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n537), .A2(KEYINPUT105), .A3(new_n571), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT105), .B1(new_n537), .B2(new_n571), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n644), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n714), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n219), .B1(new_n722), .B2(new_n467), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT106), .B1(new_n707), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n715), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n699), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n537), .A2(new_n571), .A3(KEYINPUT105), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n699), .B2(new_n719), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n467), .B(new_n713), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G29gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n706), .A4(new_n703), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n724), .A2(new_n735), .ZN(G1328gat));
  NAND3_X1  g535(.A1(new_n696), .A2(new_n220), .A3(new_n420), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT46), .Z(new_n738));
  AND2_X1   g537(.A1(new_n722), .A2(new_n420), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n220), .ZN(G1329gat));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n542), .B(new_n713), .C1(new_n729), .C2(new_n731), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(G43gat), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n696), .A2(new_n744), .A3(new_n685), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n741), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g546(.A(KEYINPUT47), .B(new_n745), .C1(new_n742), .C2(G43gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n544), .B(new_n713), .C1(new_n729), .C2(new_n731), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n696), .A2(new_n516), .A3(new_n544), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n753), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT48), .B(new_n755), .C1(new_n751), .C2(G50gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n756), .ZN(G1331gat));
  AOI21_X1  g556(.A(new_n266), .B1(new_n727), .B2(new_n728), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n657), .A2(new_n659), .A3(new_n666), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n666), .B1(new_n657), .B2(new_n659), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n645), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n671), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g564(.A(new_n420), .B(KEYINPUT107), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n763), .B2(new_n543), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n575), .A3(new_n685), .A4(new_n762), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n521), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT108), .B(G78gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n607), .A2(new_n266), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n699), .A2(new_n719), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(KEYINPUT51), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(KEYINPUT51), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n786), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n699), .A2(new_n719), .A3(new_n782), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n761), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n467), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n782), .A2(new_n668), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n671), .B(new_n792), .C1(new_n718), .C2(new_n721), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(G85gat), .B2(new_n793), .ZN(G1336gat));
  NAND2_X1  g593(.A1(new_n787), .A2(new_n789), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n766), .A2(new_n411), .A3(new_n668), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT110), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n767), .B(new_n792), .C1(new_n718), .C2(new_n721), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n411), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n783), .A2(new_n801), .A3(KEYINPUT51), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT51), .B1(new_n783), .B2(new_n801), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n792), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n420), .B(new_n805), .C1(new_n729), .C2(new_n731), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n797), .A2(new_n804), .B1(new_n806), .B2(G92gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n800), .B1(new_n807), .B2(new_n808), .ZN(G1337gat));
  AOI21_X1  g608(.A(G99gat), .B1(new_n790), .B2(new_n685), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n543), .B(new_n792), .C1(new_n718), .C2(new_n721), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(G99gat), .B2(new_n811), .ZN(G1338gat));
  OAI211_X1 g611(.A(new_n544), .B(new_n805), .C1(new_n729), .C2(new_n731), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n521), .A2(G106gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n790), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n521), .A2(G106gat), .A3(new_n761), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n804), .A2(new_n819), .B1(new_n813), .B2(G106gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n649), .A2(new_n652), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT10), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n658), .A3(new_n654), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n664), .B1(new_n657), .B2(KEYINPUT54), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n658), .B1(new_n825), .B2(new_n654), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n666), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n829), .A2(new_n266), .A3(new_n834), .A4(new_n667), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT112), .B1(new_n249), .B2(new_n251), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n244), .A2(new_n246), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n248), .A2(new_n838), .A3(new_n235), .A4(new_n250), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n261), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n265), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n668), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n719), .B1(new_n835), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n834), .A2(new_n847), .A3(new_n667), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n841), .A2(KEYINPUT113), .A3(new_n265), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n642), .A2(new_n643), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(new_n832), .B2(new_n833), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n710), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n669), .A2(new_n712), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(KEYINPUT114), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n521), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n521), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n766), .A2(new_n671), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n685), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n270), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n378), .A2(new_n521), .A3(new_n484), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n857), .A2(new_n467), .A3(new_n868), .A4(new_n858), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n766), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n330), .A3(new_n266), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(G1340gat));
  NAND2_X1  g671(.A1(new_n332), .A2(new_n334), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n873), .A3(new_n668), .ZN(new_n874));
  INV_X1    g673(.A(new_n864), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n684), .B(new_n875), .C1(new_n861), .C2(new_n862), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n668), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT116), .B1(new_n877), .B2(G120gat), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n879), .B(new_n331), .C1(new_n876), .C2(new_n668), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n878), .B2(new_n880), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n870), .B2(new_n607), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n711), .A2(G127gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n876), .B2(new_n883), .ZN(G1342gat));
  NOR4_X1   g683(.A1(new_n869), .A2(G134gat), .A3(new_n420), .A4(new_n644), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(G134gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n876), .B2(new_n719), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT117), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n885), .B(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g690(.A(G134gat), .B1(new_n865), .B2(new_n644), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(G1343gat));
  AND2_X1   g694(.A1(new_n857), .A2(new_n858), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n542), .A2(new_n521), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n467), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G141gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n700), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n898), .A2(new_n766), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n901), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n854), .ZN(new_n907));
  INV_X1    g706(.A(new_n852), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n761), .B2(new_n842), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n668), .A2(new_n843), .A3(KEYINPUT118), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n832), .A2(new_n833), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT55), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n827), .A2(new_n828), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT119), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n270), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n759), .B1(new_n916), .B2(KEYINPUT55), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n908), .B1(new_n920), .B2(new_n719), .ZN(new_n921));
  INV_X1    g720(.A(new_n607), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n521), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n875), .A2(new_n542), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n857), .A2(new_n927), .A3(new_n544), .A4(new_n858), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n926), .A2(new_n700), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n906), .B1(new_n899), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT58), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n903), .A2(new_n905), .B1(new_n904), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n266), .A3(new_n928), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n930), .A2(new_n931), .B1(new_n932), .B2(new_n934), .ZN(G1344gat));
  NOR2_X1   g734(.A1(new_n898), .A2(new_n766), .ZN(new_n936));
  INV_X1    g735(.A(G148gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n668), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n857), .A2(new_n544), .A3(new_n858), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT57), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n921), .A2(new_n922), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n645), .A2(new_n700), .A3(new_n668), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n927), .B(new_n544), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n941), .A2(new_n944), .A3(new_n668), .A4(new_n925), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n939), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n924), .A2(new_n668), .A3(new_n928), .A4(new_n925), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(new_n939), .A3(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n938), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g750(.A(KEYINPUT122), .B(new_n938), .C1(new_n946), .C2(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1345gat));
  AOI21_X1  g752(.A(G155gat), .B1(new_n936), .B2(new_n607), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n926), .A2(new_n711), .A3(new_n928), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(G155gat), .B2(new_n955), .ZN(G1346gat));
  AND3_X1   g755(.A1(new_n926), .A2(new_n719), .A3(new_n928), .ZN(new_n957));
  INV_X1    g756(.A(G162gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n719), .A2(new_n958), .A3(new_n674), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n957), .A2(new_n958), .B1(new_n898), .B2(new_n959), .ZN(G1347gat));
  NOR2_X1   g759(.A1(new_n767), .A2(new_n467), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n896), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(new_n867), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n283), .A3(new_n266), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n674), .A2(new_n467), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT124), .Z(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI211_X1 g767(.A(new_n684), .B(new_n968), .C1(new_n861), .C2(new_n862), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n700), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G169gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n965), .A2(new_n971), .ZN(G1348gat));
  AOI21_X1  g771(.A(G176gat), .B1(new_n963), .B2(new_n668), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n761), .A2(new_n299), .A3(new_n300), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n969), .B2(new_n974), .ZN(G1349gat));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n963), .A2(new_n314), .A3(new_n607), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n969), .A2(new_n711), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n976), .B(new_n977), .C1(new_n978), .C2(new_n291), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n291), .B1(new_n969), .B2(new_n711), .ZN(new_n980));
  INV_X1    g779(.A(new_n977), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT60), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n963), .A2(new_n292), .A3(new_n719), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n719), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(G190gat), .ZN(new_n987));
  AOI211_X1 g786(.A(KEYINPUT61), .B(new_n292), .C1(new_n969), .C2(new_n719), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(G1351gat));
  INV_X1    g788(.A(new_n962), .ZN(new_n990));
  INV_X1    g789(.A(G197gat), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n990), .A2(new_n991), .A3(new_n266), .A4(new_n897), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n941), .A2(new_n944), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(new_n543), .A3(new_n967), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n994), .A2(new_n700), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n995), .B2(new_n991), .ZN(G1352gat));
  NAND4_X1  g795(.A1(new_n990), .A2(new_n663), .A3(new_n668), .A4(new_n897), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  AND4_X1   g798(.A1(new_n543), .A2(new_n993), .A3(new_n668), .A4(new_n967), .ZN(new_n1000));
  OAI211_X1 g799(.A(new_n998), .B(new_n999), .C1(new_n1000), .C2(new_n663), .ZN(G1353gat));
  NAND4_X1  g800(.A1(new_n993), .A2(new_n543), .A3(new_n607), .A4(new_n967), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G211gat), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1003), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n990), .A2(new_n383), .A3(new_n607), .A4(new_n897), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(G211gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(G1354gat));
  NAND2_X1  g811(.A1(new_n719), .A2(G218gat), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT127), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n990), .A2(new_n719), .A3(new_n897), .ZN(new_n1015));
  AOI22_X1  g814(.A1(new_n994), .A2(new_n1014), .B1(new_n384), .B2(new_n1015), .ZN(G1355gat));
endmodule


