//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n213), .B(new_n219), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n217), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n202), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n208), .A2(new_n261), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n265), .A2(G150), .B1(new_n204), .B2(G20), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n254), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n201), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n253), .B1(new_n207), .B2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(new_n201), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT76), .A3(KEYINPUT9), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n267), .A2(new_n275), .ZN(new_n278));
  OR2_X1    g0078(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT77), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT66), .B1(new_n285), .B2(new_n217), .ZN(new_n286));
  AND2_X1   g0086(.A1(G1), .A2(G13), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n286), .A2(new_n290), .A3(new_n292), .A4(G274), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n286), .A2(new_n290), .ZN(new_n295));
  INV_X1    g0095(.A(G226), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n295), .A2(new_n296), .A3(new_n292), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n261), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1698), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G222), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(G223), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G77), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n302), .B(new_n304), .C1(new_n305), .C2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT67), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n285), .A2(new_n217), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n306), .B2(new_n307), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n294), .B(new_n297), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT74), .B(G200), .Z(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n316), .B2(new_n312), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n318));
  NAND3_X1  g0118(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n281), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n284), .A2(new_n317), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n282), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n312), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n276), .C1(G169), .C2(new_n312), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n286), .A2(new_n290), .A3(G244), .A4(new_n291), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT70), .B1(new_n293), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n301), .A2(G232), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n303), .A2(G238), .A3(G1698), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT71), .B(G107), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n333), .C1(new_n303), .C2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n309), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n293), .A2(new_n330), .A3(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n270), .A2(G77), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G77), .B2(new_n273), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n264), .A2(KEYINPUT72), .ZN(new_n346));
  INV_X1    g0146(.A(new_n255), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n264), .A2(KEYINPUT72), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n254), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT73), .B(new_n254), .C1(new_n345), .C2(new_n349), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n342), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n327), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n340), .B(new_n354), .C1(new_n355), .C2(new_n338), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n338), .A2(new_n316), .ZN(new_n357));
  INV_X1    g0157(.A(new_n342), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n350), .A2(new_n351), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n350), .A2(new_n351), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT75), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n315), .B1(new_n336), .B2(new_n337), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT75), .B1(new_n364), .B2(new_n354), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n336), .A2(G190), .A3(new_n337), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n323), .A2(new_n329), .A3(new_n356), .A4(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n286), .A2(new_n290), .A3(G238), .A4(new_n291), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G226), .A2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n236), .B2(G1698), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n373), .B2(new_n303), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n369), .B(new_n293), .C1(new_n374), .C2(new_n310), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n236), .A2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G226), .B2(G1698), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n370), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n309), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n369), .A4(new_n293), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT14), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(G169), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT80), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n339), .B1(new_n376), .B2(new_n385), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT80), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n286), .A2(G274), .A3(new_n290), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n292), .B1(new_n382), .B2(new_n309), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n384), .A4(new_n369), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n375), .B2(KEYINPUT13), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n396), .A2(new_n376), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n386), .A2(G169), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n399), .A2(G179), .B1(new_n400), .B2(KEYINPUT14), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT12), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n271), .B2(new_n203), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n270), .A2(KEYINPUT12), .A3(G68), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n405), .B1(new_n274), .B2(new_n203), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n264), .A2(new_n201), .B1(new_n208), .B2(G68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n208), .A2(G33), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n305), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n253), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT11), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n410), .A2(new_n411), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n406), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n396), .A2(new_n398), .A3(G190), .A4(new_n376), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n386), .A2(G200), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n414), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n299), .A2(new_n208), .A3(new_n300), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n299), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n300), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n203), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G58), .A2(G68), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT81), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(G58), .A3(G68), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n430), .A3(new_n214), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G20), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n265), .A2(G159), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n421), .B1(new_n426), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT7), .B1(new_n381), .B2(new_n208), .ZN(new_n436));
  INV_X1    g0236(.A(new_n425), .ZN(new_n437));
  OAI21_X1  g0237(.A(G68), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n431), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(KEYINPUT16), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n440), .A3(new_n253), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n259), .A2(new_n270), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n273), .B2(new_n259), .ZN(new_n443));
  INV_X1    g0243(.A(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(G223), .B(new_n444), .C1(new_n379), .C2(new_n380), .ZN(new_n445));
  OAI211_X1 g0245(.A(G226), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G87), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n448), .A2(new_n309), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n286), .A2(new_n290), .A3(G232), .A4(new_n291), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n293), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(G169), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n293), .A2(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n309), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n355), .A3(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n441), .A2(new_n443), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT18), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(G190), .A3(new_n454), .ZN(new_n458));
  OAI21_X1  g0258(.A(G200), .B1(new_n449), .B2(new_n451), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n441), .A2(new_n443), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT17), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n449), .A2(new_n313), .A3(new_n451), .ZN(new_n463));
  INV_X1    g0263(.A(G200), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n453), .B2(new_n454), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(KEYINPUT17), .A3(new_n441), .A4(new_n443), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n462), .A2(new_n467), .A3(KEYINPUT82), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT82), .B1(new_n462), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n457), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n368), .A2(new_n420), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT87), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n207), .A2(G45), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n295), .A2(new_n224), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n394), .A2(KEYINPUT85), .A3(new_n476), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT85), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n286), .A2(G274), .A3(new_n290), .ZN(new_n480));
  INV_X1    g0280(.A(new_n476), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n477), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G33), .A3(G283), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G250), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n444), .C1(new_n379), .C2(new_n380), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT4), .B1(new_n301), .B2(G244), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n309), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n483), .A2(G190), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n436), .B2(new_n437), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n264), .A2(new_n305), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT6), .ZN(new_n503));
  AND2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n502), .B1(new_n508), .B2(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n254), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n270), .A2(G97), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n207), .A2(G33), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n254), .A2(new_n270), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(new_n223), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT83), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n502), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n518));
  XNOR2_X1  g0318(.A(G97), .B(G107), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n503), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(new_n208), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n334), .B1(new_n424), .B2(new_n425), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n253), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  INV_X1    g0324(.A(new_n515), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n495), .A2(new_n516), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT86), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n528), .B(new_n464), .C1(new_n483), .C2(new_n494), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n478), .A2(new_n482), .ZN(new_n530));
  INV_X1    g0330(.A(new_n477), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n494), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT86), .B1(new_n532), .B2(G200), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n527), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  AND4_X1   g0334(.A1(new_n355), .A2(new_n530), .A3(new_n494), .A4(new_n531), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n339), .B1(new_n483), .B2(new_n494), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n535), .A2(new_n536), .B1(new_n510), .B2(new_n515), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n472), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n532), .A2(G200), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n528), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n510), .A2(KEYINPUT83), .A3(new_n515), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n532), .A2(KEYINPUT86), .A3(G200), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(new_n544), .A3(new_n545), .A4(new_n495), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT87), .A3(new_n537), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n295), .A2(new_n476), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n550));
  OAI211_X1 g0350(.A(G250), .B(new_n444), .C1(new_n379), .C2(new_n380), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G294), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n549), .A2(G264), .B1(new_n553), .B2(new_n309), .ZN(new_n554));
  AOI21_X1  g0354(.A(G169), .B1(new_n530), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n530), .A2(new_n554), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n324), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT88), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n334), .B2(G20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n496), .A2(G20), .ZN(new_n561));
  INV_X1    g0361(.A(G116), .ZN(new_n562));
  OAI22_X1  g0362(.A1(KEYINPUT23), .A2(new_n561), .B1(new_n408), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n558), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT23), .B1(new_n500), .B2(new_n208), .ZN(new_n565));
  INV_X1    g0365(.A(new_n561), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n559), .B1(new_n262), .B2(G116), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n303), .A2(new_n208), .A3(G87), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n570), .B(KEYINPUT22), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT24), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n254), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n566), .A2(new_n269), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT25), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n254), .A2(new_n270), .A3(new_n513), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(G107), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n557), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n530), .A2(new_n554), .A3(new_n313), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n556), .B2(G200), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n574), .B1(new_n569), .B2(new_n571), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n253), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n587), .A3(new_n580), .ZN(new_n588));
  OAI211_X1 g0388(.A(G238), .B(new_n444), .C1(new_n379), .C2(new_n380), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n261), .C2(new_n562), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n309), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n286), .A2(new_n290), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n473), .A2(new_n222), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n473), .A2(G274), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n316), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n497), .A2(new_n499), .A3(new_n221), .A4(new_n223), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n208), .B1(new_n370), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n408), .B2(new_n223), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n303), .A2(new_n208), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n603), .C1(new_n203), .C2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(new_n253), .B1(new_n271), .B2(new_n343), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n579), .A2(G87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n592), .A2(new_n596), .A3(G190), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n598), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n253), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n271), .A2(new_n343), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n579), .A2(new_n344), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n597), .A2(new_n339), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n592), .A2(new_n596), .A3(new_n327), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n582), .A2(new_n588), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n252), .A2(new_n217), .B1(G20), .B2(new_n562), .ZN(new_n620));
  INV_X1    g0420(.A(new_n488), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n208), .B1(new_n223), .B2(G33), .ZN(new_n622));
  OAI211_X1 g0422(.A(KEYINPUT20), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n485), .B2(new_n487), .ZN(new_n625));
  INV_X1    g0425(.A(new_n620), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n270), .A2(G116), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n579), .B2(G116), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n593), .A2(G270), .A3(new_n481), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n303), .A2(G264), .A3(G1698), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n303), .A2(G257), .A3(new_n444), .ZN(new_n634));
  INV_X1    g0434(.A(G303), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n303), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n309), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n530), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n631), .B1(new_n638), .B2(G200), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n313), .B2(new_n638), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n324), .B1(new_n636), .B2(new_n309), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n631), .A2(new_n641), .A3(new_n530), .A4(new_n632), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n339), .B1(new_n628), .B2(new_n630), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n638), .A2(new_n643), .A3(new_n644), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n640), .B(new_n642), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n619), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n471), .A2(new_n548), .A3(new_n648), .ZN(G372));
  XOR2_X1   g0449(.A(new_n616), .B(KEYINPUT89), .Z(new_n650));
  NAND4_X1  g0450(.A1(new_n546), .A2(new_n537), .A3(new_n588), .A4(new_n618), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n530), .A2(new_n554), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n339), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n530), .A2(new_n554), .A3(new_n324), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n587), .B2(new_n580), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n642), .B1(new_n646), .B2(new_n645), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n650), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n537), .A2(new_n617), .A3(new_n660), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n535), .A2(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n516), .A2(new_n526), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(KEYINPUT90), .C1(new_n535), .C2(new_n536), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n618), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n661), .B1(new_n667), .B2(new_n660), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n471), .B1(new_n659), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n329), .ZN(new_n670));
  INV_X1    g0470(.A(new_n416), .ZN(new_n671));
  INV_X1    g0471(.A(new_n419), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n356), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n468), .A2(new_n469), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n457), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n670), .B1(new_n676), .B2(new_n323), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(new_n657), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n269), .A2(new_n208), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT27), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n680), .B2(KEYINPUT27), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(G213), .B1(new_n680), .B2(KEYINPUT27), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n631), .ZN(new_n689));
  MUX2_X1   g0489(.A(new_n679), .B(new_n647), .S(new_n689), .Z(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT92), .Z(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n582), .A2(new_n588), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n587), .A2(new_n580), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n688), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n582), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n679), .A2(new_n688), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n695), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n701), .B(new_n703), .C1(new_n582), .C2(new_n688), .ZN(G399));
  INV_X1    g0504(.A(new_n211), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n599), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n215), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n548), .A2(new_n648), .A3(new_n698), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n592), .A2(new_n632), .A3(new_n596), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n530), .A3(new_n641), .A4(new_n554), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n716), .B2(new_n532), .ZN(new_n717));
  INV_X1    g0517(.A(new_n641), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n592), .A2(new_n632), .A3(new_n596), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n532), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT30), .A4(new_n556), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n355), .B1(new_n592), .B2(new_n596), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n532), .A2(new_n638), .A3(new_n652), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n717), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n688), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n713), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n688), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(KEYINPUT93), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n712), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n698), .B1(new_n659), .B2(new_n668), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n664), .A2(KEYINPUT26), .A3(new_n618), .A4(new_n666), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n660), .B1(new_n537), .B2(new_n617), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT29), .B(new_n698), .C1(new_n742), .C2(new_n659), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n711), .B1(new_n746), .B2(G1), .ZN(G364));
  NOR2_X1   g0547(.A1(new_n268), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n207), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n706), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n693), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n691), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n211), .A2(new_n303), .ZN(new_n754));
  INV_X1    g0554(.A(G355), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n755), .B1(G116), .B2(new_n211), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n705), .A2(new_n303), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G45), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n216), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n250), .A2(G45), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT95), .ZN(new_n765));
  OAI21_X1  g0565(.A(G20), .B1(new_n765), .B2(G169), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n339), .A2(KEYINPUT95), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n287), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT96), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n762), .B2(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n751), .B1(new_n764), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n327), .A2(new_n208), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n313), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G322), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n208), .A2(G190), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n355), .A2(new_n464), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G311), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n303), .B1(new_n789), .B2(G329), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n782), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n778), .A2(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G190), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n316), .A2(new_n324), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT99), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n797), .A2(new_n208), .A3(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G283), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n792), .A2(new_n313), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n787), .A2(G190), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n802), .A2(G326), .B1(G294), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n800), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n797), .A2(new_n208), .A3(new_n313), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT101), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n806), .B1(new_n801), .B2(new_n805), .C1(new_n635), .C2(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT102), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT102), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n780), .B(KEYINPUT97), .Z(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(G58), .B1(new_n798), .B2(G107), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n784), .B(KEYINPUT98), .Z(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G77), .B1(G50), .B2(new_n802), .ZN(new_n818));
  INV_X1    g0618(.A(new_n804), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n303), .B1(new_n819), .B2(new_n223), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n789), .A2(G159), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G68), .C2(new_n793), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n807), .A2(G87), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n815), .A2(new_n818), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n811), .A2(new_n812), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n777), .B1(new_n826), .B2(new_n771), .ZN(new_n827));
  INV_X1    g0627(.A(new_n774), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n691), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n753), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NOR2_X1   g0631(.A1(new_n356), .A2(new_n688), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n354), .A2(new_n688), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n367), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n832), .B1(new_n834), .B2(new_n356), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n737), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n698), .B(new_n835), .C1(new_n659), .C2(new_n668), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n751), .B1(new_n736), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n736), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n808), .A2(G107), .ZN(new_n842));
  INV_X1    g0642(.A(new_n798), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n221), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n303), .B1(new_n789), .B2(G311), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n223), .B2(new_n819), .C1(new_n780), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G283), .B2(new_n793), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n817), .A2(G116), .B1(G303), .B2(new_n802), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n842), .A2(new_n845), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n798), .A2(G68), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n303), .B1(new_n788), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n854), .A2(KEYINPUT104), .B1(G58), .B2(new_n804), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n817), .A2(G159), .B1(G150), .B2(new_n793), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n814), .A2(G143), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n802), .A2(G137), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n857), .B1(new_n861), .B2(new_n862), .C1(new_n201), .C2(new_n809), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n771), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n771), .A2(new_n772), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n751), .B1(new_n868), .B2(G77), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT103), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n866), .B(new_n870), .C1(new_n773), .C2(new_n835), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n841), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n748), .A2(new_n207), .ZN(new_n874));
  INV_X1    g0674(.A(new_n456), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT108), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n441), .A2(new_n443), .ZN(new_n877));
  INV_X1    g0677(.A(new_n686), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g0679(.A(KEYINPUT108), .B(new_n686), .C1(new_n441), .C2(new_n443), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n875), .B(new_n460), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT109), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n686), .B1(new_n441), .B2(new_n443), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(new_n876), .ZN(new_n884));
  INV_X1    g0684(.A(new_n460), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n456), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT109), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n884), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n882), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n879), .A2(new_n880), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT18), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n456), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n462), .A2(new_n467), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT106), .B1(new_n426), .B2(new_n434), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n438), .A2(new_n902), .A3(new_n439), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n903), .A3(new_n421), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n426), .A2(new_n434), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n254), .B1(new_n905), .B2(KEYINPUT16), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT107), .B1(new_n907), .B2(new_n443), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT107), .ZN(new_n909));
  INV_X1    g0709(.A(new_n443), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(new_n904), .C2(new_n906), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n452), .A2(new_n686), .A3(new_n455), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n885), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n900), .B1(new_n914), .B2(new_n888), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n878), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n470), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n899), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n712), .A2(new_n731), .A3(new_n732), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n393), .A2(new_n401), .A3(new_n419), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n698), .A2(new_n414), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n924), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n396), .A2(new_n398), .A3(G179), .A4(new_n376), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n387), .B2(new_n390), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n389), .B2(new_n392), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n419), .B(new_n926), .C1(new_n929), .C2(new_n414), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n416), .A2(new_n922), .A3(new_n419), .A4(new_n926), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n931), .A2(new_n835), .A3(new_n932), .ZN(new_n933));
  AND4_X1   g0733(.A1(KEYINPUT40), .A2(new_n920), .A3(new_n921), .A4(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n915), .B2(new_n918), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n933), .B(new_n921), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT110), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT110), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n934), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n471), .A2(new_n921), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n945), .A2(G330), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n832), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n838), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n931), .A2(new_n932), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n935), .A2(new_n936), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n894), .B2(new_n686), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT38), .B1(new_n891), .B2(new_n896), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n935), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n915), .A2(new_n918), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n898), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n671), .A2(new_n698), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n956), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n471), .A2(new_n743), .A3(new_n739), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n677), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n968), .B(new_n970), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n874), .B1(new_n948), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n971), .B2(new_n948), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n974), .A2(new_n975), .A3(G116), .A4(new_n218), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT36), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n216), .A2(G77), .A3(new_n430), .A4(new_n428), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(G50), .B2(new_n203), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(G1), .A3(new_n268), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n973), .A2(new_n977), .A3(new_n980), .ZN(G367));
  OAI21_X1  g0781(.A(new_n703), .B1(new_n582), .B2(new_n688), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n546), .B(new_n537), .C1(new_n544), .C2(new_n698), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n662), .A2(new_n698), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT44), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n982), .A2(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n701), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n692), .A2(KEYINPUT112), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n703), .B1(new_n700), .B2(new_n702), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n745), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n706), .B(KEYINPUT41), .Z(new_n997));
  OAI21_X1  g0797(.A(new_n749), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n606), .A2(new_n607), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n688), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n650), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n618), .A2(new_n1000), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1001), .A2(KEYINPUT111), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT111), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT43), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(KEYINPUT43), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n986), .A2(new_n703), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT42), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n538), .B1(new_n985), .B2(new_n656), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n688), .B2(new_n1010), .ZN(new_n1011));
  MUX2_X1   g0811(.A(new_n1005), .B(new_n1007), .S(new_n1011), .Z(new_n1012));
  NOR2_X1   g0812(.A1(new_n701), .A2(new_n986), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n998), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n381), .B1(new_n789), .B2(G137), .ZN(new_n1016));
  INV_X1    g0816(.A(G150), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n203), .B2(new_n819), .C1(new_n780), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n817), .B2(G50), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G143), .A2(new_n802), .B1(new_n793), .B2(G159), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n807), .A2(G58), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n798), .A2(G77), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n807), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1024), .A2(KEYINPUT46), .A3(new_n562), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n808), .A2(G116), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(KEYINPUT46), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT113), .B(G317), .Z(new_n1028));
  OAI221_X1 g0828(.A(new_n381), .B1(new_n1028), .B2(new_n788), .C1(new_n819), .C2(new_n334), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n817), .B2(G283), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n814), .A2(G303), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G294), .A2(new_n793), .B1(new_n802), .B2(G311), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n798), .A2(G97), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1027), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT47), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n771), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n751), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n757), .A2(new_n242), .B1(new_n705), .B2(new_n344), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n775), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n828), .C2(new_n1006), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1015), .A2(new_n1043), .ZN(G387));
  INV_X1    g0844(.A(new_n995), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n745), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n707), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n746), .B2(new_n995), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n995), .A2(new_n750), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n754), .A2(new_n708), .B1(G107), .B2(new_n211), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n758), .B1(new_n239), .B2(G45), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n708), .B(new_n759), .C1(new_n203), .C2(new_n305), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n255), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1051), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n775), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n751), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n819), .A2(new_n343), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n303), .B1(new_n1017), .B2(new_n788), .C1(new_n784), .C2(new_n203), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G50), .C2(new_n781), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G159), .A2(new_n802), .B1(new_n793), .B2(new_n260), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n807), .A2(G77), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1064), .A2(new_n1033), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n817), .A2(G303), .B1(G311), .B2(new_n793), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n802), .A2(G322), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n813), .C2(new_n1028), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(G283), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1024), .A2(new_n847), .B1(new_n1073), .B2(new_n819), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n303), .B1(new_n789), .B2(G326), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n562), .C2(new_n843), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT49), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1067), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1061), .B1(new_n1080), .B2(new_n771), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n700), .B2(new_n828), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1048), .A2(new_n1050), .A3(new_n1082), .ZN(G393));
  AOI21_X1  g0883(.A(new_n707), .B1(new_n1046), .B2(new_n992), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1046), .B2(new_n992), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n992), .A2(new_n750), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1060), .B1(G97), .B2(new_n705), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n247), .A2(new_n757), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1040), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n303), .B1(new_n789), .B2(G322), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n1024), .B2(new_n1073), .C1(new_n496), .C2(new_n843), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT116), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n784), .A2(new_n847), .B1(new_n562), .B2(new_n819), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n802), .A2(G317), .B1(new_n781), .B2(G311), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT52), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G303), .C2(new_n793), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n819), .A2(new_n305), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n381), .B(new_n1097), .C1(G143), .C2(new_n789), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n793), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n201), .C1(new_n816), .C2(new_n255), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1100), .B(new_n844), .C1(G68), .C2(new_n807), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n802), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  AOI22_X1  g0903(.A1(new_n1092), .A2(new_n1096), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n771), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1089), .B1(new_n828), .B2(new_n985), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1085), .A2(new_n1086), .A3(new_n1106), .ZN(G390));
  AOI22_X1  g0907(.A1(new_n959), .A2(new_n962), .B1(new_n953), .B2(new_n965), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n933), .A2(G330), .A3(new_n734), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n965), .B1(new_n935), .B2(new_n958), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n834), .A2(new_n356), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n698), .B(new_n1111), .C1(new_n742), .C2(new_n659), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n951), .B1(new_n1112), .B2(new_n949), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT117), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n953), .A2(new_n965), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n963), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n966), .B1(new_n899), .B2(new_n919), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n949), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n952), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1118), .A2(new_n1120), .B1(new_n735), .B2(new_n933), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT117), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n921), .A2(G330), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1126), .A2(new_n836), .A3(new_n951), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1115), .A2(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n750), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n751), .B1(new_n868), .B2(new_n260), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n852), .B1(new_n847), .B2(new_n788), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n809), .A2(new_n221), .B1(KEYINPUT119), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n817), .A2(G97), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n303), .B(new_n1097), .C1(new_n781), .C2(G116), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G283), .A2(new_n802), .B1(new_n793), .B2(new_n500), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n807), .A2(G150), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n817), .A2(new_n1141), .B1(G137), .B2(new_n793), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n804), .A2(G159), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n381), .B1(new_n789), .B2(G125), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n780), .C2(new_n853), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G128), .B2(new_n802), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1142), .B(new_n1146), .C1(new_n201), .C2(new_n843), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1132), .A2(new_n1137), .B1(new_n1139), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1130), .B1(new_n1148), .B2(new_n771), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n964), .B2(new_n773), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1129), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT120), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n471), .A2(G330), .A3(new_n921), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n969), .A2(new_n1153), .A3(new_n677), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n952), .B1(new_n735), .B2(new_n835), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n950), .B1(new_n1155), .B2(new_n1127), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n951), .B1(new_n1126), .B2(new_n836), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1157), .A2(new_n949), .A3(new_n1112), .A4(new_n1109), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1154), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1115), .A2(new_n1123), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1161));
  AND4_X1   g0961(.A1(KEYINPUT118), .A2(new_n1160), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT118), .B1(new_n1128), .B2(new_n1159), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n706), .B1(new_n1159), .B2(new_n1128), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1152), .A2(new_n1164), .ZN(G378));
  XNOR2_X1  g0965(.A(new_n1154), .B(KEYINPUT122), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT123), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n323), .A2(new_n329), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n276), .A2(new_n878), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n943), .B2(G330), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n920), .A2(KEYINPUT40), .A3(new_n921), .A4(new_n933), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n941), .B1(new_n937), .B2(new_n938), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(G330), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1171), .B(new_n1172), .Z(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n968), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n940), .A2(new_n942), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1183), .A2(G330), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n968), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1168), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1168), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1167), .B(KEYINPUT57), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT124), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1167), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n707), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1185), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT123), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1188), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT124), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT57), .A4(new_n1167), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1191), .A2(new_n1195), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1192), .A2(new_n750), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n751), .B1(new_n868), .B2(G50), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n303), .A2(G41), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT121), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1066), .B1(new_n843), .B2(new_n202), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1205), .B1(new_n1073), .B2(new_n788), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G68), .B2(new_n804), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n496), .B2(new_n780), .C1(new_n343), .C2(new_n784), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n802), .A2(G116), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1099), .B2(new_n223), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1209), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1208), .B1(new_n1215), .B2(KEYINPUT58), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n785), .A2(G137), .B1(G150), .B2(new_n804), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n781), .A2(G128), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n793), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n802), .A2(G125), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n1024), .C2(new_n1140), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n798), .A2(G159), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1216), .B1(KEYINPUT58), .B2(new_n1215), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1204), .B1(new_n1228), .B2(new_n771), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1173), .B2(new_n773), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1203), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1202), .A2(new_n1231), .ZN(G375));
  AOI21_X1  g1032(.A(new_n749), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n951), .A2(new_n772), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n751), .B1(new_n868), .B2(G68), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n808), .A2(G159), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n819), .A2(new_n201), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n381), .B(new_n1237), .C1(G128), .C2(new_n789), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n802), .A2(G132), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n1017), .C2(new_n784), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n793), .B2(new_n1141), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n814), .A2(G137), .B1(new_n798), .B2(G58), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1236), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1062), .B1(G303), .B2(new_n789), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1073), .B2(new_n780), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n817), .B2(new_n500), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G116), .A2(new_n793), .B1(new_n802), .B2(G294), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(new_n809), .C2(new_n223), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1022), .A2(new_n381), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT125), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1243), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1235), .B1(new_n1251), .B2(new_n771), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1233), .B1(new_n1234), .B2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1159), .A2(new_n997), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1156), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1254), .B2(new_n1256), .ZN(G381));
  NOR3_X1   g1057(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT126), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1202), .A2(new_n1231), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1151), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1164), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(G390), .A2(G387), .A3(G381), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .A4(new_n1264), .ZN(G407));
  NAND2_X1  g1065(.A1(new_n687), .A2(G213), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1260), .A2(new_n1263), .A3(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(G407), .A2(G213), .A3(new_n1268), .ZN(G409));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1202), .A2(G378), .A3(new_n1231), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1199), .A2(new_n750), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n1230), .C1(new_n997), .C2(new_n1193), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1263), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1266), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1159), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n707), .B1(new_n1278), .B2(new_n1256), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1256), .B2(new_n1278), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1253), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(new_n872), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n872), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1270), .B1(new_n1276), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(G387), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1287), .A2(G390), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(G390), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(G393), .B(new_n830), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1285), .A2(G2897), .A3(new_n1267), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1267), .A2(G2897), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1283), .A2(new_n1284), .A3(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1267), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1285), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1286), .A2(new_n1294), .A3(new_n1299), .A4(new_n1302), .ZN(new_n1303));
  XOR2_X1   g1103(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1304));
  AND3_X1   g1104(.A1(new_n1300), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1300), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1305), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1303), .B1(new_n1311), .B2(new_n1294), .ZN(G405));
  NOR2_X1   g1112(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1271), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1301), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1313), .A2(new_n1314), .A3(new_n1301), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1316), .A2(new_n1317), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1294), .A3(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(G402));
endmodule


