//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G143), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  OAI21_X1  g009(.A(G128), .B1(new_n189), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(G146), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n196), .B(KEYINPUT67), .C1(new_n200), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n202), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n190), .B2(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT67), .B1(new_n206), .B2(new_n196), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n194), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .B1(new_n212), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n214), .B(new_n215), .C1(KEYINPUT11), .C2(new_n213), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n212), .A2(G137), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n212), .A2(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(KEYINPUT68), .B(new_n194), .C1(new_n204), .C2(new_n207), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n210), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n210), .A2(KEYINPUT69), .A3(new_n220), .A4(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n191), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT0), .B(G128), .Z(new_n227));
  NAND2_X1  g041(.A1(new_n206), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n214), .B1(KEYINPUT11), .B2(new_n213), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n216), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(G116), .B(G119), .Z(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT2), .B(G113), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n224), .A2(new_n225), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n208), .B1(new_n241), .B2(new_n220), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n220), .A2(new_n241), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n234), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n238), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n187), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT28), .B1(new_n239), .B2(new_n222), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  INV_X1    g063(.A(G953), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G210), .ZN(new_n251));
  XOR2_X1   g065(.A(new_n251), .B(KEYINPUT27), .Z(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n252), .B(new_n253), .Z(new_n254));
  AOI21_X1  g068(.A(KEYINPUT29), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n235), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n224), .A2(new_n225), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n238), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n244), .B2(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n240), .ZN(new_n262));
  INV_X1    g076(.A(new_n254), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(KEYINPUT72), .A3(new_n263), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n255), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n240), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n224), .A2(KEYINPUT74), .A3(new_n225), .A4(new_n239), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n224), .A2(new_n225), .A3(new_n234), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n238), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n247), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n281));
  OAI21_X1  g095(.A(G472), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n258), .A2(new_n260), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n240), .A2(new_n254), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n261), .A2(KEYINPUT70), .A3(new_n240), .A4(new_n254), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n263), .B1(new_n246), .B2(new_n247), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n261), .A2(new_n292), .A3(new_n240), .A4(new_n254), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n284), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n291), .A2(new_n293), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n289), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(KEYINPUT71), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n283), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  AOI211_X1 g116(.A(KEYINPUT32), .B(new_n302), .C1(new_n295), .C2(new_n298), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n282), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  XNOR2_X1  g121(.A(G110), .B(G140), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT82), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n250), .A2(G227), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n309), .B(new_n310), .Z(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n197), .A2(new_n199), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n201), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n192), .B1(new_n315), .B2(KEYINPUT1), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n194), .B1(new_n316), .B2(new_n191), .ZN(new_n317));
  INV_X1    g131(.A(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G107), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(G107), .ZN(new_n321));
  OAI21_X1  g135(.A(G101), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(new_n318), .B2(G107), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  INV_X1    g138(.A(G107), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G104), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n323), .A2(new_n326), .A3(new_n327), .A4(new_n319), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n317), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT84), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G128), .B1(new_n200), .B2(new_n195), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n314), .A2(new_n201), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n189), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n329), .B1(new_n336), .B2(new_n194), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT84), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n313), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n210), .A2(KEYINPUT10), .A3(new_n221), .A4(new_n330), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n323), .A2(new_n326), .A3(new_n319), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(G101), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(G101), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n345), .A2(new_n342), .A3(KEYINPUT4), .A4(new_n328), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n230), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n339), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n233), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT85), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT85), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n351), .A3(new_n233), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n233), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n339), .A2(new_n354), .A3(new_n340), .A4(new_n347), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n312), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n333), .A2(new_n338), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n208), .A2(new_n330), .ZN(new_n358));
  OAI211_X1 g172(.A(KEYINPUT12), .B(new_n233), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT12), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n331), .A2(new_n332), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n337), .A2(KEYINPUT84), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n363), .B2(new_n354), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n312), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n359), .B2(new_n364), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n306), .B(new_n307), .C1(new_n356), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(new_n364), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n312), .B1(new_n372), .B2(new_n355), .ZN(new_n373));
  INV_X1    g187(.A(new_n368), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n353), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G469), .B1(new_n375), .B2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G221), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT81), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n380), .B2(new_n307), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n250), .A2(G224), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n229), .A2(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT87), .ZN(new_n388));
  INV_X1    g202(.A(G125), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(new_n194), .C1(new_n204), .C2(new_n207), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n229), .A2(new_n391), .A3(G125), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT7), .B(new_n386), .C1(new_n393), .C2(KEYINPUT88), .ZN(new_n394));
  INV_X1    g208(.A(new_n392), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n229), .B2(G125), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n397), .A2(new_n398), .A3(new_n390), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n402));
  INV_X1    g216(.A(G119), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G116), .ZN(new_n404));
  OAI211_X1 g218(.A(G113), .B(new_n404), .C1(new_n236), .C2(new_n402), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n236), .B2(new_n237), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(new_n329), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G122), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT8), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n406), .A2(new_n329), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n346), .A2(new_n238), .A3(new_n344), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n408), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT89), .A3(new_n307), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n394), .B2(new_n400), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(KEYINPUT6), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n421), .B(new_n422), .Z(new_n423));
  XOR2_X1   g237(.A(new_n393), .B(new_n386), .Z(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n401), .B2(new_n415), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n430), .A2(KEYINPUT89), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n427), .A3(new_n420), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n385), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n190), .A2(new_n434), .A3(G128), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n192), .A2(G143), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n314), .B2(new_n192), .ZN(new_n437));
  OAI211_X1 g251(.A(G134), .B(new_n435), .C1(new_n437), .C2(new_n434), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G122), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT94), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n325), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n441), .A2(new_n325), .ZN(new_n444));
  OAI221_X1 g258(.A(new_n438), .B1(G134), .B2(new_n437), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT95), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n442), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n437), .B(G134), .ZN(new_n448));
  INV_X1    g262(.A(G116), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT14), .A3(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n439), .ZN(new_n451));
  OAI211_X1 g265(.A(G107), .B(new_n450), .C1(new_n451), .C2(KEYINPUT14), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n445), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n380), .A2(G217), .A3(new_n250), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n307), .ZN(new_n459));
  INV_X1    g273(.A(G478), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT15), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT91), .B(G104), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n463), .B(new_n464), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n249), .A2(new_n250), .A3(G214), .ZN(new_n467));
  MUX2_X1   g281(.A(G143), .B(new_n190), .S(new_n467), .Z(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G125), .B(G140), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT90), .B1(new_n471), .B2(new_n201), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n201), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n468), .B(G131), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT17), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(KEYINPUT16), .ZN(new_n478));
  OR3_X1    g292(.A1(new_n389), .A2(KEYINPUT16), .A3(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n201), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n468), .A2(KEYINPUT17), .A3(G131), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(G146), .A3(new_n479), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n466), .B(new_n475), .C1(new_n477), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n471), .B(KEYINPUT19), .Z(new_n486));
  OAI211_X1 g300(.A(new_n476), .B(new_n483), .C1(G146), .C2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n487), .A2(new_n475), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n488), .B2(new_n466), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(KEYINPUT92), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT20), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n477), .A2(new_n484), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n466), .B1(new_n497), .B2(new_n475), .ZN(new_n498));
  INV_X1    g312(.A(new_n485), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n307), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT93), .B(G475), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n462), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n250), .A2(G952), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(G237), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n307), .B(new_n250), .C1(G234), .C2(G237), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n433), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT96), .B1(new_n383), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n427), .B1(new_n431), .B2(new_n420), .ZN(new_n513));
  AND4_X1   g327(.A1(new_n427), .A2(new_n417), .A3(new_n420), .A4(new_n425), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n384), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n381), .B1(new_n371), .B2(new_n376), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n504), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n296), .A2(KEYINPUT71), .A3(new_n297), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT71), .B1(new_n296), .B2(new_n297), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n300), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT32), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n299), .A2(new_n283), .A3(new_n300), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n282), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n471), .A2(new_n201), .ZN(new_n530));
  OR3_X1    g344(.A1(new_n403), .A2(KEYINPUT76), .A3(G128), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT76), .B1(new_n403), .B2(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n403), .A2(G128), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT24), .B(G110), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT77), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n403), .A2(G128), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n533), .B(new_n537), .C1(new_n538), .C2(KEYINPUT23), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n536), .B1(G110), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT77), .B1(new_n534), .B2(new_n535), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n483), .B(new_n530), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n481), .A2(new_n483), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(G110), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(new_n535), .C2(new_n534), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT22), .B(G137), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n250), .A2(G221), .A3(G234), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n547), .B(new_n548), .Z(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n545), .A3(new_n549), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n307), .ZN(new_n554));
  NOR2_X1   g368(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n555), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G217), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(G234), .B2(new_n307), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(G902), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT80), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n305), .A2(new_n521), .A3(new_n529), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  OAI21_X1  g385(.A(new_n307), .B1(new_n522), .B2(new_n523), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(new_n524), .A3(new_n569), .A4(new_n517), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT97), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n575), .A2(KEYINPUT97), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n458), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n456), .A2(KEYINPUT97), .A3(new_n575), .A4(new_n457), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n460), .A2(G902), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n580), .A2(new_n581), .B1(new_n460), .B2(new_n459), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n496), .A2(new_n502), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n516), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT34), .B(G104), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G6));
  AOI21_X1  g402(.A(G902), .B1(new_n456), .B2(new_n457), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(new_n461), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n503), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n516), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n574), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT98), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G107), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G9));
  NOR2_X1   g410(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n546), .B(new_n597), .Z(new_n598));
  INV_X1    g412(.A(new_n564), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n559), .B2(new_n561), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n573), .A2(new_n524), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n520), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT37), .B(G110), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G12));
  NOR2_X1   g420(.A1(new_n383), .A2(new_n601), .ZN(new_n607));
  INV_X1    g421(.A(new_n433), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n583), .A2(new_n462), .ZN(new_n609));
  INV_X1    g423(.A(G900), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n507), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n506), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n305), .A2(new_n529), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G128), .ZN(G30));
  NAND2_X1  g432(.A1(new_n429), .A2(new_n432), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT38), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n583), .A2(new_n590), .A3(new_n385), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(new_n601), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n613), .B(KEYINPUT39), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n517), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n620), .B(new_n622), .C1(new_n624), .C2(KEYINPUT40), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(KEYINPUT40), .B2(new_n624), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n288), .A2(new_n289), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n271), .A2(new_n272), .B1(new_n238), .B2(new_n274), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT99), .B1(new_n628), .B2(new_n254), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n254), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n307), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n527), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n314), .ZN(G45));
  NOR3_X1   g450(.A1(new_n582), .A2(new_n583), .A3(new_n614), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(KEYINPUT100), .A3(new_n433), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n584), .A2(new_n613), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n639), .B1(new_n640), .B2(new_n608), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n607), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n305), .A2(new_n529), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  AND3_X1   g458(.A1(new_n348), .A2(new_n351), .A3(new_n233), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n351), .B1(new_n348), .B2(new_n233), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n355), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n369), .A2(new_n368), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n647), .A2(new_n311), .B1(new_n648), .B2(new_n366), .ZN(new_n649));
  OAI21_X1  g463(.A(G469), .B1(new_n649), .B2(G902), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n382), .A3(new_n371), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n650), .A2(new_n371), .A3(KEYINPUT101), .A4(new_n382), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n585), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n305), .A2(new_n529), .A3(new_n569), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT41), .B(G113), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G15));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n592), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n305), .A2(new_n529), .A3(new_n569), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  NAND2_X1  g476(.A1(new_n602), .A2(new_n504), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n655), .A2(new_n515), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n305), .A2(new_n664), .A3(new_n529), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G119), .ZN(G21));
  NAND2_X1  g480(.A1(new_n462), .A2(new_n503), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n655), .A2(new_n515), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n297), .B1(new_n277), .B2(new_n254), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT102), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n297), .C1(new_n277), .C2(new_n254), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n293), .A3(new_n672), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n673), .A2(new_n300), .B1(new_n572), .B2(G472), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n668), .A2(new_n569), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  NAND4_X1  g490(.A1(new_n653), .A2(new_n433), .A3(new_n637), .A4(new_n654), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n678), .A3(new_n602), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n672), .A2(new_n293), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n628), .A2(new_n187), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n263), .B1(new_n681), .B2(new_n247), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n671), .B1(new_n682), .B2(new_n297), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n300), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n573), .A2(new_n684), .A3(new_n602), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT103), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n677), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n389), .ZN(G27));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n619), .B2(new_n385), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT104), .A4(new_n384), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n517), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n640), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n305), .A2(new_n529), .A3(new_n569), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n692), .A2(new_n640), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n304), .A2(new_n695), .A3(new_n569), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G131), .ZN(G33));
  NOR2_X1   g513(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n528), .B1(new_n527), .B2(new_n282), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n692), .A2(new_n609), .A3(new_n614), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n569), .A4(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n305), .A2(new_n529), .A3(new_n569), .A4(new_n704), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  INV_X1    g523(.A(new_n582), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n583), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n602), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n524), .B2(new_n573), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  OR3_X1    g530(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT44), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n375), .A2(KEYINPUT45), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n375), .A2(KEYINPUT45), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(G469), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(G469), .A2(G902), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT46), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n649), .A2(G469), .A3(G902), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n720), .A2(KEYINPUT46), .A3(new_n721), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n381), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(new_n623), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n690), .A2(new_n691), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n715), .B2(KEYINPUT44), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n716), .B1(new_n715), .B2(KEYINPUT44), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n717), .A2(new_n727), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G137), .ZN(G39));
  NOR4_X1   g546(.A1(new_n702), .A2(new_n569), .A3(new_n640), .A4(new_n728), .ZN(new_n733));
  NOR2_X1   g547(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n726), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G140), .ZN(G42));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n713), .A2(new_n506), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n569), .A3(new_n674), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n655), .A2(new_n384), .A3(new_n620), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT50), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT50), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n650), .A2(new_n371), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n737), .B1(new_n381), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n728), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n742), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n745), .B(new_n746), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n655), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n741), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n678), .A2(new_n573), .A3(new_n684), .A4(new_n602), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n678), .B1(new_n674), .B2(new_n602), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n750), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n527), .A2(new_n569), .A3(new_n506), .A4(new_n633), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n760), .A2(new_n761), .A3(KEYINPUT113), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT113), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n583), .A3(new_n582), .A4(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n758), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n740), .B1(new_n752), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n584), .A3(new_n763), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n655), .A2(new_n608), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n505), .B1(new_n742), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n568), .B1(new_n527), .B2(new_n282), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n754), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n766), .A2(new_n771), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n752), .A2(new_n740), .A3(new_n765), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n695), .B1(new_n756), .B2(new_n755), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n602), .A2(new_n504), .A3(new_n613), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n692), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n305), .A2(new_n529), .A3(new_n784), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n697), .A2(new_n694), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n657), .A2(new_n661), .A3(new_n665), .A4(new_n675), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n604), .A2(new_n586), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n583), .B2(new_n462), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n503), .A2(new_n590), .A3(KEYINPUT108), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT109), .B1(new_n792), .B2(new_n516), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(KEYINPUT109), .A3(new_n516), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n574), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n788), .A2(new_n570), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n708), .A2(new_n786), .A3(new_n787), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n305), .A2(new_n529), .A3(new_n616), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(new_n687), .ZN(new_n801));
  INV_X1    g615(.A(new_n677), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n756), .B2(new_n755), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n617), .A3(KEYINPUT110), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n377), .A2(new_n382), .A3(new_n601), .A4(new_n613), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT111), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n621), .A2(new_n619), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n634), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n643), .A2(KEYINPUT52), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n801), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n803), .A2(new_n617), .A3(new_n643), .A4(new_n808), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n798), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n811), .B(new_n812), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n786), .A2(new_n796), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n657), .A2(new_n661), .A3(new_n665), .A4(new_n675), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n705), .B2(new_n707), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n811), .B(KEYINPUT52), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n816), .B1(new_n825), .B2(new_n797), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n814), .A2(new_n819), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n781), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(G952), .A2(G953), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n382), .A2(new_n384), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n620), .A2(new_n568), .A3(new_n711), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n747), .A2(KEYINPUT49), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n747), .A2(KEYINPUT49), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n830), .A2(new_n831), .B1(new_n634), .B2(new_n836), .ZN(G75));
  AOI21_X1  g651(.A(new_n307), .B1(new_n826), .B2(new_n827), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n838), .B2(G210), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n423), .B(new_n424), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT55), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n839), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n250), .A2(G952), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT117), .Z(new_n844));
  AND2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(G51));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n720), .B(KEYINPUT119), .Z(new_n847));
  AND2_X1   g661(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n721), .B(KEYINPUT57), .Z(new_n849));
  NAND2_X1  g663(.A1(new_n826), .A2(new_n827), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n826), .A2(new_n827), .A3(new_n852), .A4(new_n828), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT54), .B1(new_n822), .B2(new_n816), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n855), .B2(new_n827), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n849), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n649), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n848), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n846), .B1(new_n859), .B2(new_n843), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n853), .A3(new_n851), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n649), .B1(new_n862), .B2(new_n849), .ZN(new_n863));
  OAI221_X1 g677(.A(KEYINPUT120), .B1(G952), .B2(new_n250), .C1(new_n863), .C2(new_n848), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(G54));
  AND3_X1   g679(.A1(new_n838), .A2(KEYINPUT58), .A3(G475), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n489), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n489), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(new_n868), .A3(new_n843), .ZN(G60));
  XNOR2_X1  g683(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n870));
  NAND2_X1  g684(.A1(G478), .A2(G902), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n578), .B2(new_n579), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT122), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n824), .B2(new_n829), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n844), .B1(new_n876), .B2(new_n580), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n877), .ZN(G63));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n560), .A2(new_n307), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n850), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n553), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n884), .B(new_n844), .C1(new_n598), .C2(new_n882), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT61), .Z(G66));
  AND2_X1   g700(.A1(new_n787), .A2(new_n796), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(G953), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT124), .ZN(new_n889));
  INV_X1    g703(.A(G224), .ZN(new_n890));
  OAI21_X1  g704(.A(G953), .B1(new_n508), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(G898), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n423), .B1(new_n893), .B2(G953), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n892), .B(new_n894), .Z(G69));
  AOI21_X1  g709(.A(new_n250), .B1(G227), .B2(G900), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n727), .A2(new_n773), .A3(new_n807), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n698), .A2(new_n731), .A3(new_n738), .A4(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n801), .A2(new_n643), .A3(new_n804), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n250), .A3(new_n708), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n244), .A2(new_n256), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n258), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT125), .Z(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(new_n486), .Z(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(G900), .B2(G953), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n896), .B1(new_n906), .B2(KEYINPUT127), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n899), .A2(new_n635), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT62), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n909), .B2(KEYINPUT62), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(KEYINPUT62), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n792), .A2(new_n584), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n915), .A2(new_n624), .A3(new_n728), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n702), .A2(new_n569), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n731), .A2(new_n738), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n913), .A2(new_n914), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n250), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n904), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n921), .B2(new_n906), .ZN(new_n922));
  INV_X1    g736(.A(new_n906), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n923), .B(new_n907), .C1(new_n920), .C2(new_n904), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(G72));
  NAND2_X1  g739(.A1(new_n262), .A2(new_n254), .ZN(new_n926));
  INV_X1    g740(.A(new_n887), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT63), .Z(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n898), .A2(new_n708), .A3(new_n899), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n932), .B2(new_n927), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n262), .A2(new_n254), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n843), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n627), .A2(new_n266), .A3(new_n267), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n823), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n931), .A2(new_n938), .ZN(G57));
endmodule


