//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923;
  XNOR2_X1  g000(.A(KEYINPUT68), .B(G71gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G99gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G15gat), .B(G43gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT24), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT24), .A3(new_n214), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT25), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n213), .A2(new_n215), .A3(new_n219), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(KEYINPUT25), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT66), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT27), .B(G183gat), .Z(new_n229));
  OAI21_X1  g028(.A(KEYINPUT28), .B1(new_n229), .B2(G190gat), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n216), .A2(KEYINPUT65), .A3(KEYINPUT27), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT27), .B1(new_n216), .B2(KEYINPUT65), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n217), .A4(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n225), .B(new_n226), .C1(new_n209), .C2(new_n210), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n228), .A2(new_n230), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G127gat), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n238), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n242), .A2(new_n240), .A3(KEYINPUT1), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n237), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n248), .A3(new_n236), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n207), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n205), .B1(new_n250), .B2(KEYINPUT33), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT69), .A3(KEYINPUT34), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n205), .C1(new_n250), .C2(KEYINPUT33), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT32), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n247), .A2(new_n207), .A3(new_n249), .ZN(new_n258));
  OR2_X1    g057(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n258), .B(new_n259), .C1(new_n250), .C2(new_n256), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n252), .A2(new_n262), .A3(new_n261), .A4(new_n254), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n267));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT70), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT22), .ZN(new_n271));
  INV_X1    g070(.A(G211gat), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(KEYINPUT71), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n278), .A2(new_n283), .A3(new_n279), .A4(new_n275), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G162gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G141gat), .B(G148gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(KEYINPUT2), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT76), .B(G155gat), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G162gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n291), .B2(KEYINPUT2), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n286), .B(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n293), .B1(new_n292), .B2(new_n295), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n285), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n289), .C1(new_n296), .C2(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n282), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n284), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT81), .B(new_n298), .C1(new_n285), .C2(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n277), .A2(new_n312), .A3(new_n280), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(new_n282), .C1(new_n312), .C2(new_n277), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n303), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n310), .B1(new_n315), .B2(new_n298), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n307), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G78gat), .B(G106gat), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G22gat), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT31), .B(G50gat), .Z(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n311), .A2(new_n317), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n266), .A2(new_n267), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n267), .B1(new_n266), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT35), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n301), .A2(new_n246), .A3(new_n304), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n289), .B(new_n248), .C1(new_n296), .C2(new_n297), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n334));
  AND2_X1   g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n298), .A2(new_n246), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n335), .B1(new_n340), .B2(new_n333), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(KEYINPUT5), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n333), .A2(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n332), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  INV_X1    g154(.A(new_n353), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n342), .A2(new_n356), .A3(new_n347), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(KEYINPUT6), .A3(new_n353), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n361), .B(KEYINPUT72), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n237), .A2(KEYINPUT73), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n224), .A2(new_n365), .A3(new_n236), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT29), .B(new_n362), .C1(new_n224), .C2(new_n236), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n306), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n224), .B2(new_n236), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(new_n282), .A3(new_n366), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n363), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(new_n306), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n373), .A2(new_n377), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT30), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n373), .A2(new_n377), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n360), .A2(new_n378), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n329), .A2(new_n330), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n348), .A2(KEYINPUT84), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n342), .A2(new_n388), .A3(new_n347), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n353), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n357), .A2(new_n355), .ZN(new_n391));
  INV_X1    g190(.A(new_n354), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n381), .A2(new_n378), .A3(new_n384), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n266), .A2(new_n326), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT35), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n386), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT40), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n331), .A2(new_n345), .A3(new_n343), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT39), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n335), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n356), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT83), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n406), .A3(new_n356), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n401), .A2(new_n335), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n340), .A2(new_n333), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n409), .B(KEYINPUT39), .C1(new_n410), .C2(new_n335), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n400), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n403), .A2(new_n406), .A3(new_n356), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n406), .B1(new_n403), .B2(new_n356), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n400), .B(new_n411), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n394), .B(new_n390), .C1(new_n412), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n377), .B1(new_n373), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n418), .B2(new_n373), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n379), .B1(new_n420), .B2(KEYINPUT38), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n372), .A2(new_n306), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n367), .A2(new_n368), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(KEYINPUT37), .C1(new_n306), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n373), .A2(new_n418), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n376), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n417), .A2(new_n326), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n326), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n385), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n266), .B(KEYINPUT36), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n399), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G229gat), .A2(G233gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT13), .ZN(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G22gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT91), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n439), .A2(G1gat), .ZN(new_n440));
  INV_X1    g239(.A(G8gat), .ZN(new_n441));
  INV_X1    g240(.A(G1gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n440), .B2(new_n444), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(G29gat), .A2(G36gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT14), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G29gat), .A2(G36gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT87), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(G29gat), .A3(G36gat), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n451), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G50gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G43gat), .ZN(new_n463));
  INV_X1    g262(.A(G43gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G50gat), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT15), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(new_n458), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n448), .A2(KEYINPUT88), .A3(new_n449), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n451), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n463), .A2(new_n465), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT89), .A4(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT15), .B1(new_n463), .B2(new_n465), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n466), .A2(new_n479), .A3(new_n468), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT89), .B1(new_n480), .B2(new_n473), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n467), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT15), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n476), .A2(new_n459), .A3(new_n486), .ZN(new_n487));
  NOR4_X1   g286(.A1(new_n470), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT88), .B1(new_n448), .B2(new_n449), .ZN(new_n489));
  INV_X1    g288(.A(new_n451), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n485), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n477), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT90), .A3(new_n467), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n447), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n445), .A2(new_n446), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n484), .A3(new_n494), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n437), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n436), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n482), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n495), .B2(new_n502), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT92), .B1(new_n504), .B2(new_n497), .ZN(new_n505));
  AOI221_X4 g304(.A(new_n483), .B1(new_n461), .B2(new_n466), .C1(new_n492), .C2(new_n477), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT90), .B1(new_n493), .B2(new_n467), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n503), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT92), .A4(new_n497), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n501), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n499), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n497), .A3(new_n509), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n510), .ZN(new_n519));
  AND4_X1   g318(.A1(new_n515), .A2(new_n519), .A3(KEYINPUT18), .A4(new_n501), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n500), .B1(new_n518), .B2(new_n510), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n515), .B1(new_n521), .B2(KEYINPUT18), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n514), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524));
  INV_X1    g323(.A(G197gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT11), .B(G169gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT12), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n514), .B(new_n529), .C1(new_n520), .C2(new_n522), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT94), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT94), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n523), .A2(new_n534), .A3(new_n530), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G71gat), .B(G78gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(G183gat), .B1(new_n447), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n497), .B(new_n216), .C1(new_n544), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n544), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT97), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n546), .A3(new_n547), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n557), .B2(new_n558), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT98), .B(G211gat), .Z(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n561), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n561), .B2(new_n562), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT99), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580));
  OAI211_X1 g379(.A(KEYINPUT99), .B(new_n580), .C1(new_n572), .C2(new_n573), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G99gat), .B(G106gat), .Z(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n504), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n495), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n571), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G230gat), .ZN(new_n608));
  INV_X1    g407(.A(G233gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n586), .B(new_n542), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n588), .A2(KEYINPUT10), .A3(new_n542), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n611), .A2(new_n608), .A3(new_n609), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OR3_X1    g418(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n435), .A2(new_n537), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n360), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n442), .ZN(G1324gat));
  INV_X1    g425(.A(new_n394), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n629));
  OR2_X1    g428(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n633), .B(new_n634), .C1(new_n441), .C2(new_n628), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n624), .B2(new_n433), .ZN(new_n636));
  INV_X1    g435(.A(new_n266), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n637), .A2(G15gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n624), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT101), .Z(G1326gat));
  INV_X1    g439(.A(new_n431), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n434), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n429), .A2(KEYINPUT102), .A3(new_n432), .A4(new_n433), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT103), .B1(new_n386), .B2(new_n398), .ZN(new_n650));
  INV_X1    g449(.A(new_n328), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n266), .A2(new_n326), .A3(new_n267), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n653), .A2(KEYINPUT35), .A3(new_n360), .A4(new_n627), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n390), .A2(new_n391), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n392), .A2(KEYINPUT6), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n627), .A2(new_n657), .A3(new_n397), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n330), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n646), .B1(new_n662), .B2(new_n606), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n606), .B1(new_n399), .B2(new_n434), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT44), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n536), .A2(new_n571), .A3(new_n622), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n645), .B1(new_n668), .B2(new_n360), .ZN(new_n669));
  INV_X1    g468(.A(new_n360), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n666), .A2(KEYINPUT104), .A3(new_n670), .A4(new_n667), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(G29gat), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n664), .A2(new_n667), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(G29gat), .A3(new_n360), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT45), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(G1328gat));
  OAI21_X1  g475(.A(G36gat), .B1(new_n668), .B2(new_n627), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n673), .A2(G36gat), .A3(new_n627), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT46), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(G1329gat));
  NOR3_X1   g479(.A1(new_n673), .A2(G43gat), .A3(new_n637), .ZN(new_n681));
  INV_X1    g480(.A(new_n433), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n682), .A3(new_n667), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n683), .B2(G43gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g484(.A(G50gat), .B1(new_n668), .B2(new_n326), .ZN(new_n686));
  INV_X1    g485(.A(new_n673), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT105), .B1(new_n641), .B2(G50gat), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n641), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(KEYINPUT48), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n690), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n666), .A2(new_n431), .A3(new_n667), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(KEYINPUT48), .B2(new_n694), .ZN(G1331gat));
  INV_X1    g494(.A(new_n622), .ZN(new_n696));
  NOR4_X1   g495(.A1(new_n662), .A2(new_n537), .A3(new_n607), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n670), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT106), .B(G57gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1332gat));
  NAND2_X1  g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n394), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  NOR2_X1   g502(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1333gat));
  INV_X1    g504(.A(new_n662), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n607), .A2(new_n537), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n622), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G71gat), .B1(new_n708), .B2(new_n433), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n637), .A2(G71gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n431), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g513(.A1(new_n648), .A2(new_n649), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n650), .A2(new_n661), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n606), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n537), .A2(new_n571), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT108), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n719), .A3(KEYINPUT51), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT51), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n696), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n572), .A3(new_n670), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n663), .A2(new_n622), .A3(new_n665), .A4(new_n719), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n360), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1336gat));
  OAI21_X1  g526(.A(G92gat), .B1(new_n725), .B2(new_n627), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n717), .A2(new_n719), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(KEYINPUT110), .A3(KEYINPUT51), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n394), .A2(new_n573), .A3(new_n622), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT109), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n728), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT52), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n728), .B(new_n739), .C1(new_n722), .C2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1337gat));
  INV_X1    g540(.A(G99gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n742), .A3(new_n266), .ZN(new_n743));
  OAI21_X1  g542(.A(G99gat), .B1(new_n725), .B2(new_n433), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1338gat));
  OAI21_X1  g544(.A(G106gat), .B1(new_n725), .B2(new_n326), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n326), .A2(new_n696), .A3(G106gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n720), .B2(new_n721), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT111), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n746), .A2(new_n752), .A3(new_n749), .A4(new_n747), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n732), .A2(new_n733), .A3(new_n748), .ZN(new_n755));
  OAI21_X1  g554(.A(G106gat), .B1(new_n725), .B2(new_n641), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT53), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n758), .ZN(G1339gat));
  NAND2_X1  g558(.A1(new_n623), .A2(new_n536), .ZN(new_n760));
  INV_X1    g559(.A(new_n528), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n436), .B1(new_n519), .B2(new_n496), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n496), .A2(new_n498), .A3(new_n437), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n532), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n619), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n615), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n613), .A2(new_n614), .A3(new_n610), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT54), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n768), .B(KEYINPUT55), .C1(new_n770), .C2(new_n615), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n620), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n770), .B2(new_n615), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n603), .A2(new_n605), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n533), .A2(new_n535), .A3(new_n774), .A4(new_n778), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n532), .A2(new_n622), .A3(new_n764), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n765), .A2(KEYINPUT113), .A3(new_n622), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n780), .B1(new_n786), .B2(new_n606), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n760), .B1(new_n787), .B2(new_n571), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n394), .A2(new_n360), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n431), .A2(new_n637), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(KEYINPUT114), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n796), .B2(new_n536), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n653), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n536), .A2(G113gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT115), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(G1340gat));
  OR3_X1    g600(.A1(new_n798), .A2(G120gat), .A3(new_n696), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n794), .A2(new_n622), .A3(new_n795), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n803), .A2(new_n804), .A3(G120gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n803), .B2(G120gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(G1341gat));
  INV_X1    g606(.A(new_n571), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n796), .A2(new_n238), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n653), .A3(new_n571), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n238), .B2(new_n810), .ZN(G1342gat));
  NOR3_X1   g610(.A1(new_n798), .A2(G134gat), .A3(new_n606), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT56), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n796), .B2(new_n606), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1343gat));
  INV_X1    g614(.A(new_n606), .ZN(new_n816));
  INV_X1    g615(.A(new_n772), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n533), .A2(new_n535), .A3(new_n778), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n818), .B2(new_n782), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n808), .B1(new_n819), .B2(new_n780), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n760), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT57), .B1(new_n821), .B2(new_n641), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  INV_X1    g622(.A(new_n326), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n788), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n789), .A2(new_n433), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G141gat), .B1(new_n827), .B2(new_n536), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n682), .A2(new_n326), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT118), .Z(new_n830));
  AND2_X1   g629(.A1(new_n790), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(G141gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n537), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT58), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n828), .B(new_n833), .C1(new_n835), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1344gat));
  INV_X1    g639(.A(G148gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n831), .A2(new_n841), .A3(new_n622), .ZN(new_n842));
  INV_X1    g641(.A(new_n827), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT59), .B(new_n841), .C1(new_n843), .C2(new_n622), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n818), .A2(new_n782), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n606), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  INV_X1    g647(.A(new_n780), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT119), .B1(new_n819), .B2(new_n780), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n808), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n760), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n641), .A2(KEYINPUT57), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n788), .A2(new_n824), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n853), .A2(new_n854), .B1(new_n855), .B2(KEYINPUT57), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n622), .A3(new_n826), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n845), .B1(new_n857), .B2(G148gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n842), .B1(new_n844), .B2(new_n858), .ZN(G1345gat));
  AOI21_X1  g658(.A(new_n290), .B1(new_n831), .B2(new_n571), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n571), .A2(new_n290), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT120), .Z(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n843), .B2(new_n862), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n831), .B2(new_n816), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n816), .A2(G162gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n843), .B2(new_n865), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n627), .A2(new_n670), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n788), .A2(new_n653), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n209), .A3(new_n537), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n788), .A2(new_n791), .A3(new_n867), .ZN(new_n870));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n536), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1348gat));
  AOI21_X1  g671(.A(G176gat), .B1(new_n868), .B2(new_n622), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT121), .Z(new_n874));
  NOR3_X1   g673(.A1(new_n870), .A2(new_n210), .A3(new_n696), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(G1349gat));
  INV_X1    g675(.A(new_n229), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n868), .A2(KEYINPUT122), .A3(new_n877), .A4(new_n571), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n788), .A2(new_n877), .A3(new_n653), .A4(new_n867), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n808), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G183gat), .B1(new_n870), .B2(new_n808), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(KEYINPUT123), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n217), .A3(new_n816), .ZN(new_n886));
  OAI21_X1  g685(.A(G190gat), .B1(new_n870), .B2(new_n606), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(KEYINPUT61), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(KEYINPUT61), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G1351gat));
  NAND2_X1  g689(.A1(new_n867), .A2(new_n433), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n856), .A2(new_n537), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n788), .A2(new_n829), .A3(new_n867), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n788), .A2(KEYINPUT124), .A3(new_n829), .A4(new_n867), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n537), .A2(new_n525), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n893), .A2(new_n525), .B1(new_n898), .B2(new_n899), .ZN(G1352gat));
  NOR3_X1   g699(.A1(new_n894), .A2(G204gat), .A3(new_n696), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT62), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n856), .A2(new_n622), .A3(new_n892), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G204gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1353gat));
  NAND2_X1  g704(.A1(new_n853), .A2(new_n854), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n855), .A2(KEYINPUT57), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n571), .A4(new_n892), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n856), .A2(KEYINPUT126), .A3(new_n571), .A4(new_n892), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(G211gat), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT63), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n910), .A2(new_n911), .A3(new_n914), .A4(G211gat), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n896), .A2(new_n272), .A3(new_n571), .A4(new_n897), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT125), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n915), .A3(new_n917), .ZN(G1354gat));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n856), .A2(new_n919), .A3(new_n892), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n856), .B2(new_n892), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n606), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n816), .A2(new_n273), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n922), .A2(new_n273), .B1(new_n898), .B2(new_n923), .ZN(G1355gat));
endmodule


