//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G210), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(G237), .A3(G953), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT26), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G101), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT28), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n193), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n199), .A2(new_n201), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G137), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT65), .B1(new_n207), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT64), .B1(new_n193), .B2(G146), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n204), .B(new_n201), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n203), .A2(new_n206), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n215), .A2(new_n218), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n210), .A2(new_n214), .A3(new_n212), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G131), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n215), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n199), .A2(new_n233), .B1(new_n235), .B2(new_n206), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT66), .B1(new_n239), .B2(G116), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(G116), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT2), .A2(G113), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT2), .A2(G113), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n244), .A2(new_n249), .A3(new_n245), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n238), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n253), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT67), .B1(new_n207), .B2(new_n219), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n225), .A2(new_n226), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .A4(new_n237), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n192), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n255), .B(new_n237), .C1(new_n207), .C2(new_n219), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(new_n192), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n191), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n238), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n256), .A2(new_n258), .A3(new_n237), .A4(KEYINPUT30), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n253), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n190), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n259), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT31), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT68), .B(new_n191), .C1(new_n260), .C2(new_n262), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n271), .A3(new_n275), .A4(new_n259), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n265), .A2(new_n273), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G472), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n271), .B1(new_n260), .B2(new_n262), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n269), .A2(new_n259), .A3(new_n191), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT29), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n256), .A2(new_n258), .A3(new_n237), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n253), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n192), .B1(new_n289), .B2(new_n259), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n262), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n285), .B2(new_n286), .ZN(new_n294));
  OAI21_X1  g108(.A(G472), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n277), .A2(KEYINPUT32), .A3(new_n278), .A4(new_n279), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(G234), .B2(new_n279), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(G953), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(G221), .A3(G234), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT22), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(G137), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n200), .B2(G119), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n239), .A2(KEYINPUT70), .A3(G128), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n307), .B(new_n308), .C1(new_n239), .C2(G128), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT24), .B(G110), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n239), .B2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n239), .A2(G128), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n311), .B1(G110), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT71), .B(G125), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n319), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT71), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G125), .A2(G140), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n322), .B(KEYINPUT16), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n319), .B2(new_n323), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n322), .B1(new_n333), .B2(KEYINPUT16), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n321), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n196), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n327), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n329), .B1(new_n337), .B2(G140), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT16), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT72), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n330), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G146), .A3(new_n321), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n318), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n196), .B(new_n320), .C1(new_n340), .C2(new_n330), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n309), .A2(new_n310), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT73), .B(G110), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(new_n314), .A3(new_n313), .A4(new_n315), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g166(.A1(G125), .A2(G140), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n332), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n332), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n196), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n305), .B1(new_n343), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n341), .B2(new_n321), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n317), .B1(new_n361), .B2(new_n344), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n342), .A2(new_n351), .A3(new_n356), .A4(new_n349), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n304), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n359), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n359), .B2(new_n364), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n300), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT77), .B(new_n300), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  INV_X1    g184(.A(new_n299), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n359), .A2(new_n279), .A3(new_n364), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(KEYINPUT25), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n359), .A2(new_n374), .A3(new_n364), .A4(new_n279), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n297), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n361), .B2(new_n344), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n336), .A2(KEYINPUT93), .A3(new_n342), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n301), .A3(G214), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n193), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n193), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n387), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n213), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  MUX2_X1   g205(.A(new_n391), .B(new_n388), .S(KEYINPUT17), .Z(new_n392));
  NAND3_X1  g206(.A1(new_n381), .A2(new_n382), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n386), .A2(new_n387), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT90), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT18), .A3(G131), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n356), .B1(new_n196), .B2(new_n333), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n399), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n393), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n396), .B1(new_n393), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n279), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT95), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(new_n279), .C1(new_n404), .C2(new_n405), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT94), .B(G475), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n396), .A3(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n388), .A2(new_n390), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n388), .B2(new_n390), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n354), .B2(new_n355), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n338), .A2(KEYINPUT19), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT92), .B1(new_n421), .B2(new_n196), .ZN(new_n422));
  AND4_X1   g236(.A1(KEYINPUT92), .A2(new_n419), .A3(new_n420), .A4(new_n196), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n342), .B(new_n417), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n403), .ZN(new_n425));
  INV_X1    g239(.A(new_n396), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n413), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT20), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n432), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G128), .B(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n193), .A2(G128), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n436), .B(G134), .C1(KEYINPUT13), .C2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G122), .ZN(new_n439));
  INV_X1    g253(.A(G107), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n209), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n435), .B(new_n209), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n242), .A2(KEYINPUT14), .A3(G122), .ZN(new_n445));
  INV_X1    g259(.A(new_n439), .ZN(new_n446));
  OAI211_X1 g260(.A(G107), .B(new_n445), .C1(new_n446), .C2(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n439), .A2(new_n440), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(new_n298), .A3(G953), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n450), .B(new_n452), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n279), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n412), .A2(new_n434), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n301), .A2(G952), .ZN(new_n459));
  NAND2_X1  g273(.A1(G234), .A2(G237), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(G902), .A3(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(G898), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT3), .B1(new_n395), .B2(G107), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n440), .A3(G104), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n395), .A2(G107), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n469), .A2(new_n471), .A3(new_n270), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n395), .A2(G107), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n440), .A2(G104), .ZN(new_n475));
  OAI21_X1  g289(.A(G101), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n252), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G113), .B1(new_n245), .B2(KEYINPUT5), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n242), .A2(G119), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n240), .B2(new_n243), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n480), .B2(KEYINPUT5), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT78), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n469), .A2(new_n471), .A3(new_n485), .A4(new_n472), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(G101), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n473), .A2(KEYINPUT4), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n487), .A2(new_n488), .B1(new_n251), .B2(new_n252), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n484), .A2(new_n490), .A3(G101), .A4(new_n486), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n482), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G122), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT82), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n487), .A2(new_n488), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n253), .A3(new_n491), .ZN(new_n498));
  INV_X1    g312(.A(new_n482), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT82), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n494), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n225), .A2(new_n337), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n199), .A2(new_n233), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n235), .A2(new_n206), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n319), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n301), .A2(G224), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n512), .B(new_n513), .Z(new_n514));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT83), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n503), .A2(new_n507), .A3(new_n517), .A4(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n244), .A2(KEYINPUT5), .A3(new_n245), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n478), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n480), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n477), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n519), .A2(new_n522), .B1(new_n249), .B2(new_n480), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n473), .A2(new_n476), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n252), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT85), .B(new_n529), .C1(new_n481), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n493), .B(KEYINPUT8), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n513), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n508), .B2(new_n511), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT7), .B1(new_n513), .B2(KEYINPUT88), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(KEYINPUT88), .B2(new_n513), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n539), .A2(KEYINPUT87), .B1(new_n512), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n536), .A2(new_n542), .A3(new_n543), .A4(new_n506), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n279), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n544), .B2(new_n279), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n516), .B(new_n518), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G210), .B1(G237), .B2(G902), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n544), .A2(new_n279), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT89), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n546), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n555), .A2(new_n550), .A3(new_n518), .A4(new_n516), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n466), .B(new_n468), .C1(new_n552), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n497), .A2(new_n236), .A3(new_n491), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n530), .A2(new_n225), .A3(KEYINPUT79), .A4(KEYINPUT10), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT79), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT10), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n207), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n230), .A2(new_n215), .ZN(new_n564));
  INV_X1    g378(.A(new_n203), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n223), .B1(new_n565), .B2(new_n199), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n530), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n558), .A2(new_n563), .A3(new_n564), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n530), .A2(new_n225), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n204), .B1(new_n221), .B2(new_n222), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n203), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n529), .B1(new_n573), .B2(new_n223), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n231), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n207), .A2(new_n529), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n579), .A2(KEYINPUT80), .A3(KEYINPUT12), .A4(new_n231), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n576), .B(new_n564), .C1(new_n567), .C2(new_n578), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT80), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n570), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G140), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n301), .A2(G227), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n587), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n558), .A2(new_n563), .A3(new_n569), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n231), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n570), .A2(KEYINPUT81), .A3(new_n589), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n588), .A2(new_n596), .A3(G469), .ZN(new_n597));
  INV_X1    g411(.A(G469), .ZN(new_n598));
  INV_X1    g412(.A(new_n581), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n582), .A2(KEYINPUT80), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n590), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n594), .B2(new_n570), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n598), .B(new_n279), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(G469), .A2(G902), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n597), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G221), .B1(new_n451), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n379), .A2(new_n458), .A3(new_n557), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NOR2_X1   g424(.A1(new_n377), .A2(new_n607), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n277), .A2(new_n279), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n611), .A2(new_n612), .A3(new_n280), .A4(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n367), .A2(new_n368), .B1(new_n373), .B2(new_n375), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n616), .A2(new_n370), .A3(new_n606), .A4(new_n605), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n280), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT96), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n452), .B2(KEYINPUT97), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n453), .B(new_n620), .Z(new_n621));
  NOR2_X1   g435(.A1(new_n455), .A2(G902), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n454), .A2(new_n455), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT98), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n454), .A2(new_n625), .A3(new_n455), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n621), .A2(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n412), .B2(new_n434), .ZN(new_n628));
  INV_X1    g442(.A(new_n466), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n468), .B1(new_n552), .B2(new_n556), .ZN(new_n630));
  AND4_X1   g444(.A1(KEYINPUT99), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT99), .B1(new_n557), .B2(new_n628), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n615), .B(new_n619), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  AOI21_X1  g449(.A(new_n457), .B1(new_n431), .B2(new_n433), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n412), .A2(new_n630), .A3(new_n629), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n615), .A3(new_n619), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n343), .A2(new_n358), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n305), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n300), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n376), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n606), .A3(new_n605), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n618), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n557), .A3(new_n458), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  AOI22_X1  g464(.A1(new_n373), .A2(new_n375), .B1(new_n643), .B2(new_n300), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n607), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n652), .A2(new_n630), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT100), .B(G900), .Z(new_n654));
  AOI21_X1  g468(.A(new_n462), .B1(new_n464), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n636), .A2(new_n412), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n636), .A2(new_n412), .A3(KEYINPUT101), .A4(new_n656), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n653), .A2(new_n297), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT102), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XOR2_X1   g477(.A(new_n655), .B(KEYINPUT39), .Z(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n607), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT105), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT105), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n667), .A2(KEYINPUT40), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n552), .A2(new_n556), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT38), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n410), .B1(new_n406), .B2(KEYINPUT95), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n677), .A2(new_n409), .B1(new_n431), .B2(new_n433), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n457), .A2(new_n468), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n676), .A2(new_n678), .A3(new_n645), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n289), .A2(new_n259), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n191), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n272), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(G902), .B1(new_n683), .B2(KEYINPUT103), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(KEYINPUT103), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n282), .A2(new_n296), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT104), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n282), .A2(new_n686), .A3(new_n689), .A4(new_n296), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n673), .A2(new_n680), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  NAND2_X1  g507(.A1(new_n412), .A2(new_n434), .ZN(new_n694));
  INV_X1    g508(.A(new_n627), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n630), .A2(new_n694), .A3(new_n695), .A4(new_n656), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n628), .A2(KEYINPUT106), .A3(new_n630), .A4(new_n656), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n297), .A2(new_n652), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  OAI21_X1  g516(.A(new_n279), .B1(new_n601), .B2(new_n602), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n606), .A3(new_n603), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n297), .A2(new_n378), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n631), .B2(new_n632), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND2_X1  g524(.A1(new_n637), .A2(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NOR2_X1   g526(.A1(new_n705), .A2(new_n651), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n557), .A2(new_n458), .A3(new_n297), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  NAND2_X1  g529(.A1(new_n278), .A2(new_n279), .ZN(new_n716));
  INV_X1    g530(.A(new_n276), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n191), .B1(new_n290), .B2(new_n262), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n273), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n717), .B1(new_n719), .B2(KEYINPUT107), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n273), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n716), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT108), .B(G472), .Z(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n277), .B2(new_n279), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n377), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n679), .B1(new_n412), .B2(new_n434), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n705), .A2(new_n466), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n727), .A2(new_n674), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  AND2_X1   g545(.A1(new_n630), .A2(new_n706), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n678), .A2(new_n627), .A3(new_n655), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n723), .A2(new_n651), .A3(new_n726), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(G125), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G27));
  NOR2_X1   g551(.A1(new_n607), .A2(KEYINPUT110), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n552), .A2(new_n467), .A3(new_n556), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n605), .B2(new_n606), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n628), .A2(new_n656), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n296), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n296), .A2(new_n746), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n282), .A3(new_n295), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n378), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n749), .B2(new_n378), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n742), .B(new_n745), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n379), .A2(new_n742), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n744), .B1(new_n754), .B2(new_n743), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n659), .A2(new_n660), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n758), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n659), .A2(new_n660), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT113), .A3(new_n379), .A4(new_n742), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(new_n606), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n588), .A2(new_n596), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n598), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT46), .B1(new_n769), .B2(new_n604), .ZN(new_n770));
  INV_X1    g584(.A(new_n603), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n604), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n765), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n665), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n678), .A2(new_n695), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n651), .B1(new_n614), .B2(new_n280), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .A4(new_n780), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n739), .B(KEYINPUT114), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n776), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  AOI211_X1 g601(.A(KEYINPUT47), .B(new_n765), .C1(new_n772), .C2(new_n773), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n743), .A2(new_n297), .A3(new_n378), .A4(new_n739), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n789), .B(new_n790), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  AND3_X1   g610(.A1(new_n297), .A2(new_n630), .A3(new_n652), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n734), .A2(new_n628), .A3(new_n656), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n761), .A2(new_n797), .B1(new_n798), .B2(new_n732), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n606), .A2(new_n651), .A3(new_n605), .A4(new_n656), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n728), .A2(new_n800), .A3(new_n674), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n691), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n701), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n701), .A2(new_n661), .A3(new_n735), .A4(new_n802), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n804), .B2(new_n806), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n753), .A2(new_n755), .B1(new_n760), .B2(new_n762), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n714), .A2(new_n730), .A3(new_n648), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n708), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n636), .A2(new_n412), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n678), .B2(new_n627), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n615), .A2(new_n619), .A3(new_n814), .A4(new_n557), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n609), .A2(new_n815), .A3(new_n711), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n412), .A2(new_n434), .A3(new_n457), .A4(new_n656), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n739), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n700), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n819), .A2(new_n818), .A3(new_n739), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n733), .A2(new_n734), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n810), .A2(new_n817), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n809), .A2(new_n827), .A3(KEYINPUT53), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n812), .A2(new_n816), .A3(new_n825), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n810), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n802), .A2(new_n661), .A3(new_n735), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n806), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n803), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n830), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n828), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n691), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n739), .A2(new_n377), .A3(new_n461), .A4(new_n705), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n678), .A3(new_n627), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n739), .A2(new_n705), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n778), .A2(new_n462), .A3(new_n779), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n734), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n778), .A2(new_n462), .A3(new_n779), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n676), .A2(new_n468), .A3(new_n706), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT50), .A4(new_n727), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n778), .A2(new_n462), .A3(new_n727), .A4(new_n779), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n848), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n846), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT47), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n774), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n704), .A2(new_n603), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n856), .A2(new_n788), .B1(new_n606), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n847), .A2(new_n859), .A3(new_n727), .A4(new_n785), .ZN(new_n860));
  INV_X1    g674(.A(new_n785), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n854), .A2(KEYINPUT51), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT51), .B1(new_n854), .B2(new_n863), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n847), .A2(new_n727), .A3(new_n732), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n459), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n840), .A2(new_n628), .A3(new_n841), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n751), .A2(new_n752), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT48), .ZN(new_n870));
  INV_X1    g684(.A(new_n844), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n867), .B(new_n868), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n864), .A2(new_n865), .A3(new_n874), .ZN(new_n875));
  AND4_X1   g689(.A1(KEYINPUT53), .A2(new_n836), .A3(new_n810), .A4(new_n831), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n809), .A2(new_n827), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n877), .B2(new_n830), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n839), .B(new_n875), .C1(new_n878), .C2(new_n829), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT119), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n378), .A2(new_n467), .A3(new_n606), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n857), .B(KEYINPUT49), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n777), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n840), .A2(new_n885), .A3(new_n676), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(G75));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n828), .A2(new_n838), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G902), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n894), .B2(new_n187), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n503), .A2(new_n507), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n514), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT55), .Z(new_n898));
  AND2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n895), .A2(new_n898), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n301), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  INV_X1    g716(.A(new_n803), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n835), .A2(KEYINPUT117), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n906), .A2(new_n830), .A3(new_n832), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n827), .B2(new_n836), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT54), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n839), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n604), .B(KEYINPUT57), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n911), .A2(new_n912), .B1(new_n602), .B2(new_n601), .ZN(new_n913));
  INV_X1    g727(.A(new_n894), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n769), .B(KEYINPUT121), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n901), .B1(new_n913), .B2(new_n916), .ZN(G54));
  NAND4_X1  g731(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .A4(new_n428), .ZN(new_n918));
  INV_X1    g732(.A(new_n901), .ZN(new_n919));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n413), .B(new_n427), .C1(new_n894), .C2(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT59), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n621), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n828), .A2(new_n829), .A3(new_n838), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n829), .B1(new_n828), .B2(new_n838), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n919), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n839), .B1(new_n878), .B2(new_n829), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n621), .B1(new_n930), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT122), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n830), .B1(new_n906), .B2(new_n832), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n829), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n924), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n621), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n901), .B1(new_n910), .B2(new_n925), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n932), .A2(new_n941), .ZN(G63));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n365), .A2(new_n366), .ZN(new_n944));
  INV_X1    g758(.A(new_n893), .ZN(new_n945));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n919), .ZN(new_n949));
  INV_X1    g763(.A(new_n643), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n945), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n943), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n951), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n919), .A4(new_n948), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(G66));
  INV_X1    g769(.A(new_n817), .ZN(new_n956));
  NAND2_X1  g770(.A1(G224), .A2(G953), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n956), .A2(G953), .B1(new_n465), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n896), .B1(G898), .B2(new_n301), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(G69));
  NAND2_X1  g774(.A1(new_n267), .A2(new_n268), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT123), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n421), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  INV_X1    g778(.A(new_n669), .ZN(new_n965));
  INV_X1    g779(.A(new_n739), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n379), .A3(new_n966), .A4(new_n814), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n795), .A2(new_n786), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n799), .A2(new_n701), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n970), .A3(new_n692), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n692), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n964), .B1(new_n974), .B2(G953), .ZN(new_n975));
  NAND2_X1  g789(.A1(G900), .A2(G953), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n795), .A2(new_n786), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n810), .A2(new_n969), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n728), .A2(new_n674), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n776), .A2(new_n979), .A3(new_n869), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n977), .B(new_n978), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n976), .B(new_n963), .C1(new_n983), .C2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n301), .B1(G227), .B2(G900), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G72));
  NAND4_X1  g801(.A1(new_n968), .A2(new_n817), .A3(new_n971), .A4(new_n973), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n191), .B1(new_n269), .B2(new_n259), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n990), .B1(new_n983), .B2(new_n956), .ZN(new_n996));
  INV_X1    g810(.A(new_n284), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n901), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n878), .ZN(new_n999));
  INV_X1    g813(.A(new_n990), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n997), .A2(new_n1000), .A3(new_n992), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n992), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n995), .A2(new_n998), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT127), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n993), .A2(new_n994), .B1(new_n999), .B2(new_n1001), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1006), .A2(new_n1007), .A3(new_n998), .A4(new_n1003), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1008), .ZN(G57));
endmodule


