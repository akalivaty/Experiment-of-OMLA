//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  AND2_X1   g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(new_n203), .C2(new_n202), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT88), .ZN(new_n211));
  AND2_X1   g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT15), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n211), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  INV_X1    g027(.A(G29gat), .ZN(new_n229));
  INV_X1    g028(.A(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n231), .A2(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(KEYINPUT88), .A3(new_n220), .A4(new_n214), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  INV_X1    g034(.A(new_n214), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n223), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n237), .A2(KEYINPUT87), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n222), .B1(new_n237), .B2(KEYINPUT87), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n235), .B1(new_n234), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n210), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT89), .B(new_n210), .C1(new_n241), .C2(new_n242), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n207), .A2(new_n248), .A3(new_n209), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n207), .B2(new_n209), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n240), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n245), .A2(new_n246), .A3(new_n247), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n234), .A2(new_n240), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n257), .A2(new_n249), .A3(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(KEYINPUT17), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n259), .A2(new_n260), .B1(new_n207), .B2(new_n209), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(KEYINPUT89), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(KEYINPUT18), .A3(new_n246), .A4(new_n245), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n249), .B2(new_n250), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n253), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n246), .B(KEYINPUT13), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT11), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT86), .ZN(new_n271));
  XNOR2_X1  g070(.A(G169gat), .B(G197gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT12), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n256), .A2(new_n263), .A3(new_n267), .A4(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT91), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  AND2_X1   g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(KEYINPUT24), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n290), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(KEYINPUT65), .A3(new_n287), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(KEYINPUT23), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n289), .A2(new_n298), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n303), .B(new_n283), .C1(new_n287), .C2(new_n286), .ZN(new_n308));
  INV_X1    g107(.A(new_n293), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(new_n292), .B2(KEYINPUT24), .ZN(new_n311));
  OR3_X1    g110(.A1(new_n292), .A2(new_n310), .A3(KEYINPUT24), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n290), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n304), .A2(new_n303), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(KEYINPUT68), .A3(new_n298), .A4(new_n289), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n307), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n283), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n286), .B1(new_n318), .B2(KEYINPUT26), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n286), .A2(KEYINPUT26), .ZN(new_n322));
  MUX2_X1   g121(.A(new_n321), .B(new_n320), .S(new_n322), .Z(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT69), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n325), .A2(new_n326), .A3(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT28), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n323), .B(new_n294), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n317), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n332), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(G127gat), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(KEYINPUT71), .B(G134gat), .C1(new_n332), .C2(KEYINPUT1), .ZN(new_n343));
  INV_X1    g142(.A(G127gat), .ZN(new_n344));
  INV_X1    g143(.A(G134gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(KEYINPUT72), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT72), .B1(new_n342), .B2(new_n347), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n317), .B(new_n330), .C1(new_n350), .C2(new_n349), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G15gat), .B(G43gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n356), .B(KEYINPUT32), .C1(new_n358), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT34), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n355), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n353), .ZN(new_n369));
  AOI211_X1 g168(.A(KEYINPUT34), .B(new_n354), .C1(new_n352), .C2(new_n355), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n363), .A3(new_n365), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT36), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(KEYINPUT73), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n371), .A2(new_n363), .A3(new_n377), .A4(new_n365), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT74), .B1(new_n366), .B2(new_n372), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n366), .A2(new_n372), .A3(KEYINPUT74), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n375), .B1(new_n386), .B2(KEYINPUT36), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT31), .B(G50gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G228gat), .ZN(new_n391));
  INV_X1    g190(.A(G233gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(G155gat), .B(G162gat), .Z(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n395), .B(KEYINPUT78), .C1(KEYINPUT2), .C2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G141gat), .ZN(new_n400));
  INV_X1    g199(.A(G141gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G148gat), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT2), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G155gat), .B(G162gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(KEYINPUT79), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G141gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n400), .B1(new_n410), .B2(new_n399), .ZN(new_n411));
  OR3_X1    g210(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n412));
  INV_X1    g211(.A(G155gat), .ZN(new_n413));
  INV_X1    g212(.A(G162gat), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n397), .A2(new_n405), .B1(new_n411), .B2(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT80), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422));
  AND2_X1   g221(.A1(G211gat), .A2(G218gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(G211gat), .A2(G218gat), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n425), .B(new_n426), .C1(KEYINPUT22), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(KEYINPUT22), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n430), .B2(KEYINPUT82), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n428), .B2(new_n429), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n422), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n421), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n430), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n435), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n422), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n394), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT3), .B1(new_n437), .B2(new_n422), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n393), .B1(new_n441), .B2(new_n420), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n390), .B1(new_n445), .B2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n439), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n416), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT80), .B1(new_n406), .B2(new_n416), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n434), .A2(new_n435), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n443), .B1(new_n453), .B2(new_n394), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n445), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n446), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(G22gat), .B1(new_n445), .B2(KEYINPUT83), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n455), .A3(new_n447), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n454), .A2(new_n455), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n390), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n342), .A2(new_n347), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n420), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n417), .A2(KEYINPUT3), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n342), .B(new_n347), .C1(new_n420), .C2(new_n435), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n344), .B1(new_n343), .B2(new_n346), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n419), .A2(new_n475), .A3(new_n421), .A4(new_n348), .ZN(new_n476));
  OAI221_X1 g275(.A(new_n469), .B1(new_n470), .B2(new_n471), .C1(new_n476), .C2(new_n468), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n417), .A2(new_n342), .A3(new_n347), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n464), .B1(new_n479), .B2(new_n467), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT81), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n477), .B(new_n482), .C1(new_n481), .C2(new_n480), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n466), .A2(KEYINPUT4), .A3(new_n420), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n471), .B2(new_n470), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n476), .A2(new_n468), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n478), .A4(new_n464), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G1gat), .B(G29gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT0), .ZN(new_n491));
  XNOR2_X1  g290(.A(G57gat), .B(G85gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT75), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n317), .B2(new_n330), .ZN(new_n497));
  INV_X1    g296(.A(G226gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n392), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n331), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n331), .A2(new_n496), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n437), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n499), .B2(new_n497), .ZN(new_n505));
  INV_X1    g304(.A(new_n437), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G64gat), .B(G92gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n504), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n504), .B2(new_n507), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n507), .A4(new_n511), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT4), .B1(new_n351), .B2(new_n451), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n465), .B1(new_n522), .B2(new_n485), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n486), .A2(new_n487), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT84), .A3(new_n465), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT39), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT85), .B1(new_n528), .B2(new_n494), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT39), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT84), .B1(new_n526), .B2(new_n465), .ZN(new_n531));
  AOI211_X1 g330(.A(new_n524), .B(new_n464), .C1(new_n486), .C2(new_n487), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT85), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(new_n493), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n479), .A2(new_n467), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n530), .B1(new_n537), .B2(new_n464), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n525), .A2(new_n527), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n521), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  AOI211_X1 g340(.A(KEYINPUT40), .B(new_n541), .C1(new_n529), .C2(new_n535), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n495), .B(new_n520), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n504), .A2(new_n544), .A3(new_n507), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n502), .A2(new_n506), .A3(new_n503), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n505), .B2(new_n437), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n545), .A2(new_n510), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n504), .A2(new_n507), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT37), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT38), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n545), .A2(new_n510), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n549), .A2(KEYINPUT38), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n483), .A2(new_n493), .A3(new_n488), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n495), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n489), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n560), .A3(new_n512), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n463), .B1(new_n543), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n559), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n563));
  INV_X1    g362(.A(new_n463), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n387), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NOR4_X1   g365(.A1(new_n379), .A2(new_n463), .A3(new_n383), .A4(new_n381), .ZN(new_n567));
  INV_X1    g366(.A(new_n563), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT35), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n373), .A3(new_n374), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n282), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575));
  AOI21_X1  g374(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G71gat), .B(G78gat), .ZN(new_n579));
  XOR2_X1   g378(.A(G57gat), .B(G64gat), .Z(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n582));
  INV_X1    g381(.A(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  XOR2_X1   g390(.A(G127gat), .B(G155gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT93), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT94), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n581), .A2(KEYINPUT95), .A3(new_n584), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT95), .B1(new_n581), .B2(new_n584), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n251), .B1(KEYINPUT21), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n589), .B(new_n590), .ZN(new_n601));
  INV_X1    g400(.A(new_n594), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n595), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n600), .B1(new_n595), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n575), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n595), .A2(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n599), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n595), .A2(new_n603), .A3(new_n600), .ZN(new_n609));
  INV_X1    g408(.A(new_n575), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT41), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT96), .Z(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G99gat), .B(G106gat), .Z(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT98), .B(G92gat), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT8), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  OAI211_X1 g425(.A(G85gat), .B(G92gat), .C1(new_n626), .C2(KEYINPUT7), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT7), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(KEYINPUT97), .A3(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n627), .A2(new_n630), .B1(new_n626), .B2(KEYINPUT7), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n619), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  INV_X1    g432(.A(new_n619), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n620), .A2(new_n621), .B1(KEYINPUT8), .B2(new_n623), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  OAI22_X1  g436(.A1(new_n257), .A2(new_n637), .B1(new_n614), .B2(new_n613), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT99), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  OAI221_X1 g439(.A(new_n640), .B1(new_n614), .B2(new_n613), .C1(new_n257), .C2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n637), .B1(new_n241), .B2(new_n242), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G190gat), .B(G218gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n618), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n618), .A4(new_n648), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G230gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n392), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n580), .A2(new_n579), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n625), .A2(new_n631), .A3(new_n619), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n585), .A2(new_n632), .A3(new_n636), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT10), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n632), .A2(new_n636), .A3(KEYINPUT10), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(new_n596), .A3(new_n597), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n658), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n663), .A2(new_n664), .A3(new_n657), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT101), .ZN(new_n673));
  XOR2_X1   g472(.A(G176gat), .B(G204gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n671), .A2(new_n676), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n612), .A2(new_n655), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n574), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n559), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT102), .B(G1gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1324gat));
  INV_X1    g485(.A(new_n683), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT103), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n687), .A2(new_n688), .A3(new_n520), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n520), .A3(new_n690), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n208), .B1(new_n687), .B2(new_n520), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n697), .B(new_n691), .C1(new_n693), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n683), .B2(new_n387), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n385), .A2(G15gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n683), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n683), .A2(new_n564), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(new_n612), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n681), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n655), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT105), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n574), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n229), .A3(new_n560), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT107), .B1(new_n569), .B2(new_n572), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n380), .A2(new_n384), .A3(new_n564), .A4(new_n382), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n571), .B1(new_n715), .B2(new_n563), .ZN(new_n716));
  INV_X1    g515(.A(new_n570), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n568), .A2(new_n717), .A3(KEYINPUT35), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n566), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT44), .B1(new_n721), .B2(new_n655), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n655), .A2(KEYINPUT44), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n566), .B2(new_n573), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n267), .ZN(new_n726));
  INV_X1    g525(.A(new_n254), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(KEYINPUT18), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(KEYINPUT91), .A3(new_n256), .A4(new_n274), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n277), .A2(new_n278), .ZN(new_n730));
  AOI221_X4 g529(.A(KEYINPUT106), .B1(new_n268), .B2(new_n275), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n276), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n707), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n559), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n713), .A2(new_n739), .ZN(G1328gat));
  INV_X1    g539(.A(new_n520), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n710), .A2(G36gat), .A3(new_n741), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n743), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(KEYINPUT108), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(KEYINPUT108), .ZN(new_n747));
  OAI221_X1 g546(.A(new_n742), .B1(new_n743), .B2(new_n744), .C1(new_n746), .C2(new_n747), .ZN(G1329gat));
  NOR4_X1   g547(.A1(new_n722), .A2(new_n387), .A3(new_n724), .A4(new_n736), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT109), .B1(new_n749), .B2(new_n215), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n711), .A2(new_n215), .A3(new_n386), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n749), .B2(new_n215), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI221_X1 g553(.A(new_n751), .B1(KEYINPUT109), .B2(KEYINPUT47), .C1(new_n749), .C2(new_n215), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1330gat));
  OAI21_X1  g555(.A(new_n216), .B1(new_n710), .B2(new_n564), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n463), .A2(G50gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n738), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1331gat));
  NOR4_X1   g560(.A1(new_n735), .A2(new_n612), .A3(new_n655), .A4(new_n680), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n721), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT111), .B1(new_n721), .B2(new_n762), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n560), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g568(.A(KEYINPUT49), .B(G64gat), .C1(new_n767), .C2(new_n520), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT49), .B(G64gat), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n765), .A2(new_n766), .A3(new_n741), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n770), .A2(new_n772), .ZN(G1333gat));
  NOR2_X1   g572(.A1(new_n385), .A2(G71gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(G71gat), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n765), .A2(new_n387), .A3(new_n766), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n775), .B(KEYINPUT50), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n463), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g583(.A1(new_n735), .A2(new_n706), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n721), .A2(new_n655), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n721), .A2(new_n788), .A3(new_n655), .A4(new_n785), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n559), .A2(G85gat), .A3(new_n680), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n681), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n722), .A2(new_n724), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n560), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(new_n621), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n741), .A2(G92gat), .A3(new_n680), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n786), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n798), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n721), .A2(new_n655), .A3(new_n785), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n797), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n722), .A2(new_n741), .A3(new_n724), .A4(new_n792), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n802), .A2(KEYINPUT113), .B1(new_n803), .B2(new_n620), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n805), .B(new_n797), .C1(new_n799), .C2(new_n801), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n789), .A3(new_n796), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n808), .B(new_n809), .C1(new_n803), .C2(new_n620), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1337gat));
  NOR3_X1   g610(.A1(new_n385), .A2(G99gat), .A3(new_n680), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n787), .A2(new_n789), .A3(new_n812), .ZN(new_n813));
  NOR4_X1   g612(.A1(new_n722), .A2(new_n387), .A3(new_n724), .A4(new_n792), .ZN(new_n814));
  INV_X1    g613(.A(G99gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT114), .ZN(G1338gat));
  NAND2_X1  g616(.A1(new_n793), .A2(new_n463), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n564), .A2(new_n680), .A3(G106gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n787), .A2(new_n789), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(G106gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n793), .B2(new_n463), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n821), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT115), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n822), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n829), .B1(new_n799), .B2(new_n801), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT53), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n828), .A3(new_n831), .ZN(G1339gat));
  AOI21_X1  g631(.A(new_n246), .B1(new_n262), .B2(new_n245), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT119), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n833), .A2(KEYINPUT119), .B1(new_n265), .B2(new_n266), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n273), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n733), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n665), .A2(new_n667), .A3(new_n658), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(KEYINPUT54), .A3(new_n668), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n842), .B(new_n658), .C1(new_n665), .C2(new_n667), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(KEYINPUT117), .A3(new_n675), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT117), .B1(new_n843), .B2(new_n675), .ZN(new_n845));
  OAI211_X1 g644(.A(KEYINPUT55), .B(new_n841), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n675), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(KEYINPUT117), .A3(new_n675), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT55), .A4(new_n841), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n855), .A2(new_n677), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n839), .A2(new_n655), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n838), .A2(new_n680), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n735), .B2(new_n859), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT120), .B(new_n861), .C1(new_n863), .C2(new_n655), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n281), .A2(KEYINPUT106), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n733), .A2(new_n732), .A3(new_n276), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n859), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n839), .A2(new_n681), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n655), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n865), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n864), .A2(new_n871), .A3(new_n612), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n866), .A2(new_n867), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n682), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n682), .A2(KEYINPUT116), .A3(new_n873), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n520), .A2(new_n559), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n570), .ZN(new_n882));
  AOI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n735), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n715), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n282), .A2(new_n337), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1340gat));
  AOI21_X1  g685(.A(G120gat), .B1(new_n882), .B2(new_n681), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n680), .A2(new_n335), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(G1341gat));
  NAND2_X1  g688(.A1(new_n882), .A2(new_n706), .ZN(new_n890));
  XOR2_X1   g689(.A(KEYINPUT71), .B(G127gat), .Z(new_n891));
  NOR2_X1   g690(.A1(new_n612), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n890), .A2(new_n891), .B1(new_n884), .B2(new_n892), .ZN(G1342gat));
  INV_X1    g692(.A(new_n881), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n895));
  INV_X1    g694(.A(new_n655), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n570), .A3(G134gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n655), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n900), .B2(G134gat), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n894), .A2(new_n897), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1343gat));
  NAND2_X1  g702(.A1(new_n387), .A2(new_n463), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n881), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n282), .A2(G141gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT58), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n387), .A2(new_n880), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n876), .A2(new_n877), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n868), .A2(new_n869), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n860), .B1(new_n911), .B2(new_n896), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n706), .B1(new_n912), .B2(KEYINPUT120), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n871), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n909), .B1(new_n914), .B2(new_n564), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n858), .B(KEYINPUT122), .Z(new_n916));
  AOI21_X1  g715(.A(new_n678), .B1(new_n847), .B2(new_n854), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n281), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n869), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n896), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n706), .B1(new_n920), .B2(new_n861), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT57), .B(new_n463), .C1(new_n910), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n908), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT123), .B1(new_n923), .B2(new_n281), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n564), .B1(new_n872), .B2(new_n878), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n925), .B2(KEYINPUT57), .ZN(new_n926));
  INV_X1    g725(.A(new_n908), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n926), .A2(KEYINPUT123), .A3(new_n281), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n410), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n907), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n410), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n923), .B2(new_n735), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n905), .A2(new_n906), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT58), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1344gat));
  OR4_X1    g734(.A1(G148gat), .A2(new_n881), .A3(new_n680), .A4(new_n904), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT59), .B(new_n399), .C1(new_n923), .C2(new_n681), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT57), .B1(new_n914), .B2(new_n564), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n682), .A2(new_n282), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n909), .B(new_n463), .C1(new_n921), .C2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n681), .A3(new_n927), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n942), .B2(G148gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n936), .B1(new_n937), .B2(new_n943), .ZN(G1345gat));
  INV_X1    g743(.A(new_n923), .ZN(new_n945));
  OAI21_X1  g744(.A(G155gat), .B1(new_n945), .B2(new_n612), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n905), .A2(new_n413), .A3(new_n706), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1346gat));
  OAI21_X1  g747(.A(G162gat), .B1(new_n945), .B2(new_n896), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n905), .A2(new_n414), .A3(new_n655), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n741), .A2(new_n560), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n879), .A2(new_n567), .A3(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n953), .A2(new_n284), .A3(new_n282), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n914), .A2(new_n560), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n741), .A2(new_n570), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(KEYINPUT125), .A3(new_n957), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n735), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n954), .B1(new_n962), .B2(new_n284), .ZN(G1348gat));
  OAI21_X1  g762(.A(G176gat), .B1(new_n953), .B2(new_n680), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n681), .A2(new_n285), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G1349gat));
  OAI21_X1  g766(.A(G183gat), .B1(new_n953), .B2(new_n612), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n612), .A2(new_n325), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n955), .A2(new_n957), .A3(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT60), .ZN(new_n972));
  AOI22_X1  g771(.A1(new_n968), .A2(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(G1350gat));
  OAI21_X1  g774(.A(G190gat), .B1(new_n953), .B2(new_n896), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n655), .A2(new_n328), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n965), .B2(new_n978), .ZN(G1351gat));
  NOR2_X1   g778(.A1(new_n904), .A2(new_n741), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n955), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n981), .A2(new_n873), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n387), .A2(new_n952), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n941), .B(new_n984), .C1(new_n925), .C2(new_n909), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n281), .A2(G197gat), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n982), .A2(G197gat), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(G1352gat));
  NOR2_X1   g787(.A1(new_n680), .A2(G204gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n955), .A2(new_n980), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g789(.A(new_n990), .B(KEYINPUT62), .Z(new_n991));
  NAND3_X1  g790(.A1(new_n939), .A2(new_n681), .A3(new_n941), .ZN(new_n992));
  OAI21_X1  g791(.A(G204gat), .B1(new_n992), .B2(new_n983), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1353gat));
  OR3_X1    g793(.A1(new_n981), .A2(G211gat), .A3(new_n612), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n985), .A2(new_n612), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n997));
  OAI211_X1 g796(.A(KEYINPUT63), .B(G211gat), .C1(new_n985), .C2(new_n612), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n995), .B1(new_n997), .B2(new_n999), .ZN(G1354gat));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n896), .B1(new_n985), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1002), .B1(new_n1001), .B2(new_n985), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G218gat), .ZN(new_n1004));
  OR3_X1    g803(.A1(new_n981), .A2(G218gat), .A3(new_n896), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1355gat));
endmodule


