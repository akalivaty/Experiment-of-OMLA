//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT71), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT72), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n461), .A2(new_n462), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G138), .A4(new_n460), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(new_n504), .B2(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n508), .B2(G62), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(G543), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n506), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT73), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n514));
  OAI211_X1 g089(.A(G62), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n501), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT74), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n505), .A2(new_n507), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n518), .A2(G88), .A3(new_n512), .A4(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n506), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n511), .A2(new_n517), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n519), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  OAI211_X1 g107(.A(KEYINPUT76), .B(G543), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(new_n512), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT75), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n508), .A2(new_n539), .A3(G63), .A4(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n508), .A2(G89), .A3(new_n519), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n535), .A2(new_n541), .A3(new_n545), .ZN(G168));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  INV_X1    g122(.A(G77), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n536), .A2(new_n547), .B1(new_n548), .B2(new_n506), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  OAI221_X1 g126(.A(new_n551), .B1(new_n548), .B2(new_n506), .C1(new_n536), .C2(new_n547), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(G651), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n530), .B2(new_n533), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n508), .A2(G90), .A3(new_n519), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n560));
  INV_X1    g135(.A(new_n533), .ZN(new_n561));
  OAI21_X1  g136(.A(G52), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT78), .B1(new_n562), .B2(new_n556), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n553), .B1(new_n559), .B2(new_n563), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  AOI22_X1  g140(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n510), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n534), .A2(G43), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n508), .A2(new_n519), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G81), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(G188));
  OAI211_X1 g152(.A(G53), .B(G543), .C1(new_n531), .C2(new_n532), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n508), .A2(G91), .A3(new_n519), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n510), .C2(new_n581), .ZN(G299));
  NAND3_X1  g157(.A1(new_n535), .A2(new_n541), .A3(new_n545), .ZN(G286));
  OAI21_X1  g158(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n508), .A2(G87), .A3(new_n519), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n523), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT79), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n584), .A2(new_n585), .A3(new_n589), .A4(new_n586), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(G288));
  OAI211_X1 g166(.A(G61), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n518), .A2(G86), .A3(new_n512), .A4(new_n519), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n523), .A2(G48), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n510), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n534), .A2(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n569), .A2(G85), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G290));
  NAND3_X1  g179(.A1(new_n508), .A2(G92), .A3(new_n519), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n508), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n560), .A2(new_n561), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n510), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT80), .B1(new_n614), .B2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  MUX2_X1   g191(.A(KEYINPUT80), .B(new_n615), .S(new_n616), .Z(G284));
  MUX2_X1   g192(.A(KEYINPUT80), .B(new_n615), .S(new_n616), .Z(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n580), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n508), .A2(G65), .ZN(new_n623));
  NAND2_X1  g198(.A1(G78), .A2(G543), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n510), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(G868), .B2(new_n626), .ZN(G297));
  OAI21_X1  g202(.A(new_n619), .B1(G868), .B2(new_n626), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n614), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n614), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT81), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(KEYINPUT81), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G868), .C2(new_n572), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g211(.A(new_n465), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n496), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n485), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n473), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n460), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(G2096), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n653), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n667), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n676), .B(new_n678), .Z(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(G166), .A2(G16), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G16), .B2(G22), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n587), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT88), .A4(new_n586), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G6), .B(G305), .S(G16), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n702), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n711), .A2(KEYINPUT34), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G24), .ZN(new_n718));
  XNOR2_X1  g293(.A(G290), .B(KEYINPUT87), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1986), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n485), .A2(G131), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(G107), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G2105), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G119), .B2(new_n473), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XOR2_X1   g307(.A(new_n731), .B(new_n732), .Z(new_n733));
  NOR3_X1   g308(.A1(new_n717), .A2(new_n721), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT34), .B1(new_n711), .B2(new_n716), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT25), .Z(new_n746));
  AOI22_X1  g321(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n460), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n485), .B2(G139), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n722), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n722), .B2(G33), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n614), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G4), .B2(G16), .ZN(new_n757));
  OAI22_X1  g332(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT30), .B(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n759), .A2(new_n722), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n646), .B2(new_n722), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n722), .A2(G32), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n485), .A2(G141), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n473), .A2(G129), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n637), .A2(G105), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n767), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n766), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n722), .A2(G26), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT28), .Z(new_n782));
  NAND3_X1  g357(.A1(new_n482), .A2(new_n484), .A3(G140), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n784));
  INV_X1    g359(.A(G116), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G2105), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G128), .B2(new_n473), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n782), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n722), .B1(KEYINPUT24), .B2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(KEYINPUT24), .B2(G34), .ZN(new_n792));
  INV_X1    g367(.A(G160), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2084), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n780), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n758), .A2(new_n765), .A3(new_n779), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n703), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n626), .B2(new_n703), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1956), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n722), .A2(G35), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n722), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT29), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n804), .B2(G2090), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT97), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT97), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n804), .A2(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n722), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n722), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n797), .A2(new_n806), .A3(new_n807), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n753), .A2(new_n754), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT93), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n703), .A2(G5), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G171), .B2(new_n703), .ZN(new_n820));
  INV_X1    g395(.A(G1961), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G168), .A2(new_n703), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n703), .B2(G21), .ZN(new_n824));
  INV_X1    g399(.A(G1966), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n826), .B(new_n827), .C1(new_n755), .C2(new_n757), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n703), .A2(G19), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n572), .B2(new_n703), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT91), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1341), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n818), .A2(new_n822), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n815), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n734), .A2(new_n737), .A3(new_n738), .A4(new_n741), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n744), .A2(new_n834), .A3(new_n835), .ZN(G150));
  INV_X1    g411(.A(G150), .ZN(G311));
  NAND2_X1  g412(.A1(new_n614), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n568), .A2(new_n570), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n534), .A2(G55), .B1(new_n569), .B2(G93), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(new_n510), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n567), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n571), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  AOI21_X1  g424(.A(G860), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n845), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT98), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT99), .ZN(G145));
  XNOR2_X1  g431(.A(new_n487), .B(new_n793), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n646), .ZN(new_n858));
  INV_X1    g433(.A(new_n788), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n774), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n768), .A2(new_n788), .A3(new_n773), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n860), .A2(G164), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(G164), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n751), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n861), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n489), .A2(new_n492), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n497), .B1(new_n480), .B2(G138), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n749), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n860), .A2(G164), .A3(new_n861), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n485), .A2(G142), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G118), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(G2105), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G130), .B2(new_n473), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n864), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n864), .B2(new_n873), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n639), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n879), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n749), .B(KEYINPUT92), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n870), .B2(new_n872), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n862), .A2(new_n863), .A3(new_n749), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n639), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n864), .A2(new_n873), .A3(new_n879), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n882), .A2(new_n890), .A3(new_n730), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT100), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n730), .B1(new_n882), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n858), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n882), .A2(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n729), .ZN(new_n897));
  INV_X1    g472(.A(new_n858), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n897), .A2(KEYINPUT100), .A3(new_n898), .A4(new_n891), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n894), .A2(new_n899), .A3(new_n895), .A4(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G395));
  XNOR2_X1  g480(.A(new_n847), .B(new_n631), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n626), .B1(new_n609), .B2(new_n613), .ZN(new_n907));
  NAND2_X1  g482(.A1(G79), .A2(G543), .ZN(new_n908));
  INV_X1    g483(.A(G66), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n536), .B2(new_n909), .ZN(new_n910));
  AOI22_X1  g485(.A1(G54), .A2(new_n534), .B1(new_n910), .B2(G651), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n607), .A2(new_n608), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(G299), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT102), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n614), .B2(G299), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n907), .A2(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n911), .A2(new_n912), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT102), .B1(new_n922), .B2(new_n626), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n921), .A2(KEYINPUT103), .A3(KEYINPUT41), .A4(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n914), .A2(new_n916), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n920), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n919), .B1(new_n930), .B2(new_n906), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  XOR2_X1   g507(.A(G303), .B(G305), .Z(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n708), .A2(G290), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n708), .A2(G290), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n934), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n935), .A3(new_n938), .ZN(new_n940));
  INV_X1    g515(.A(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT104), .B1(new_n941), .B2(new_n936), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n942), .A3(new_n933), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n932), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n932), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(G868), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n845), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(G868), .B2(new_n949), .ZN(G295));
  OAI21_X1  g525(.A(new_n948), .B1(G868), .B2(new_n949), .ZN(G331));
  NOR2_X1   g526(.A1(G301), .A2(G286), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n558), .B1(new_n555), .B2(new_n557), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n562), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G168), .B1(new_n955), .B2(new_n553), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n847), .B(KEYINPUT105), .C1(new_n952), .C2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n847), .B1(new_n952), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g533(.A1(G301), .A2(G286), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(G168), .A3(new_n553), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n846), .A3(new_n960), .A4(new_n844), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n929), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n918), .A2(new_n958), .A3(new_n961), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n944), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n895), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n944), .B1(new_n964), .B2(new_n965), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n939), .A2(new_n943), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n958), .A2(new_n961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n917), .A2(new_n925), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n920), .A2(KEYINPUT41), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n917), .B1(new_n963), .B2(new_n957), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n966), .A3(new_n978), .A4(new_n895), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n969), .A2(new_n970), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n966), .A3(new_n895), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR3_X1    g559(.A1(new_n967), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n980), .B1(new_n987), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT107), .B(G1384), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(G164), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G160), .A2(G40), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n774), .B(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n730), .A2(new_n732), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n730), .A2(new_n732), .ZN(new_n997));
  INV_X1    g572(.A(G2067), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n788), .B(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(G290), .B(G1986), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n869), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n992), .B1(new_n1007), .B2(new_n989), .ZN(new_n1008));
  INV_X1    g583(.A(new_n990), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n869), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1971), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n992), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n495), .A2(new_n498), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT50), .B(G1384), .C1(new_n1013), .C2(new_n866), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT115), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n869), .A2(new_n1016), .A3(new_n1006), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n1015), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G2090), .B1(new_n1020), .B2(KEYINPUT116), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1012), .A2(new_n1015), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1011), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1005), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n706), .A2(G1976), .A3(new_n707), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n588), .A2(new_n1028), .A3(new_n590), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1013), .B2(new_n866), .ZN(new_n1031));
  INV_X1    g606(.A(G40), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n466), .A2(new_n469), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1025), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1030), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n595), .B2(new_n598), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n510), .B1(new_n592), .B2(new_n593), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n596), .A2(new_n597), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1041), .A2(new_n1042), .A3(G1981), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1038), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n595), .A2(new_n598), .A3(new_n1039), .ZN(new_n1045));
  OAI21_X1  g620(.A(G1981), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1047), .A3(new_n1034), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT49), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(KEYINPUT111), .A3(new_n1047), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1037), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT108), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1017), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1007), .A2(KEYINPUT108), .A3(KEYINPUT50), .ZN(new_n1060));
  AOI211_X1 g635(.A(G2090), .B(new_n992), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1061), .B2(new_n1011), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT109), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1062), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1074));
  INV_X1    g649(.A(G2090), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1033), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1011), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1025), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT110), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1026), .B(new_n1056), .C1(new_n1072), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(new_n1033), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n821), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n989), .B1(G164), .B2(G1384), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(new_n1010), .A3(new_n812), .A4(new_n1033), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n466), .A2(KEYINPUT123), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n466), .A2(KEYINPUT123), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n812), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1089));
  NOR4_X1   g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n469), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n991), .A3(new_n1010), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1082), .A2(G301), .A3(new_n1086), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1031), .A2(KEYINPUT45), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1008), .A2(KEYINPUT53), .A3(new_n812), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n992), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1086), .B(new_n1094), .C1(new_n1095), .C2(G1961), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT54), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1080), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n992), .A2(G2084), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1093), .A2(new_n1083), .A3(new_n1033), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1074), .A2(new_n1104), .B1(new_n825), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1025), .B1(new_n1106), .B2(G168), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1103), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1966), .B1(new_n1008), .B2(new_n1093), .ZN(new_n1109));
  OAI21_X1  g684(.A(G286), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT51), .B(new_n1025), .C1(new_n1106), .C2(G168), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1111), .A2(KEYINPUT122), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1074), .A2(new_n1104), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1105), .A2(new_n825), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(G168), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n1110), .A3(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1107), .A2(new_n1102), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1082), .A2(new_n1086), .A3(new_n1091), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1124), .B2(G171), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1096), .A2(G171), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1099), .A2(new_n1098), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n626), .B(KEYINPUT57), .ZN(new_n1128));
  INV_X1    g703(.A(G1956), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1033), .B(new_n1057), .C1(new_n1014), .C2(KEYINPUT115), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1008), .A2(new_n1010), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1128), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1132), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n922), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1095), .A2(G1348), .B1(G2067), .B2(new_n1052), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1128), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1132), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1083), .A2(new_n1010), .A3(new_n994), .A4(new_n1033), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(G1341), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1052), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n571), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1149), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1151));
  AND2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1144), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1052), .A2(G2067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1081), .B2(new_n755), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n922), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n614), .B1(new_n1138), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1160), .A2(new_n1162), .B1(new_n1161), .B2(new_n1138), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1139), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1101), .A2(new_n1122), .A3(new_n1127), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT122), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1119), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT62), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT116), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(new_n1075), .A3(new_n1023), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1025), .B1(new_n1173), .B2(new_n1077), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1005), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1056), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1171), .A2(new_n1097), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1167), .A2(new_n1170), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1165), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(G8), .B(G168), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1056), .B(new_n1181), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1062), .A2(new_n1005), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT63), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1071), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1073), .A2(new_n1078), .A3(KEYINPUT110), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1188), .A2(new_n1189), .A3(new_n1056), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1183), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1036), .A2(new_n1030), .ZN(new_n1192));
  AOI21_X1  g767(.A(KEYINPUT111), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1193));
  AND4_X1   g768(.A1(KEYINPUT111), .A2(new_n1044), .A3(new_n1047), .A4(new_n1034), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1192), .B(new_n1035), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1191), .B1(new_n1195), .B2(new_n1180), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT118), .ZN(new_n1198));
  NOR2_X1   g773(.A1(G288), .A2(G1976), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1200), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1043), .B(KEYINPUT113), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT114), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1199), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT114), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1205), .A2(new_n1206), .A3(new_n1202), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1034), .B(KEYINPUT112), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1204), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1187), .A2(new_n1197), .A3(new_n1198), .A4(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1209), .A2(new_n1190), .A3(new_n1196), .ZN(new_n1211));
  AOI22_X1  g786(.A1(new_n1182), .A2(new_n1183), .B1(KEYINPUT63), .B2(new_n1185), .ZN(new_n1212));
  OAI21_X1  g787(.A(KEYINPUT118), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1002), .B1(new_n1179), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1000), .A2(new_n993), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT48), .ZN(new_n1217));
  INV_X1    g792(.A(new_n993), .ZN(new_n1218));
  OR3_X1    g793(.A1(new_n1218), .A2(G1986), .A3(G290), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1220), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1221));
  NOR3_X1   g796(.A1(new_n1218), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT46), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1223), .B1(new_n993), .B2(new_n994), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n999), .A2(new_n768), .A3(new_n773), .ZN(new_n1225));
  OAI22_X1  g800(.A1(new_n1222), .A2(new_n1224), .B1(new_n1225), .B2(new_n1218), .ZN(new_n1226));
  XOR2_X1   g801(.A(new_n1226), .B(KEYINPUT47), .Z(new_n1227));
  NOR2_X1   g802(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n995), .A2(new_n999), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n997), .B1(new_n1229), .B2(new_n993), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n788), .A2(G2067), .ZN(new_n1231));
  OR3_X1    g806(.A1(new_n1230), .A2(KEYINPUT125), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(KEYINPUT125), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(new_n993), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1234), .A2(KEYINPUT126), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1236));
  NAND4_X1  g811(.A1(new_n1232), .A2(new_n1236), .A3(new_n993), .A4(new_n1233), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1228), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT127), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1215), .A2(new_n1239), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g815(.A1(new_n969), .A2(new_n979), .ZN(new_n1242));
  INV_X1    g816(.A(G227), .ZN(new_n1243));
  NAND2_X1  g817(.A1(new_n1243), .A2(G319), .ZN(new_n1244));
  NOR3_X1   g818(.A1(G229), .A2(G401), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g819(.A1(new_n900), .A2(new_n1242), .A3(new_n1245), .ZN(G225));
  INV_X1    g820(.A(G225), .ZN(G308));
endmodule


