//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  OR3_X1    g002(.A1(new_n202), .A2(KEYINPUT95), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n202), .B2(KEYINPUT95), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT96), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(KEYINPUT96), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G127gat), .B(G155gat), .Z(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT100), .ZN(new_n215));
  XOR2_X1   g014(.A(G57gat), .B(G64gat), .Z(new_n216));
  XNOR2_X1  g015(.A(G71gat), .B(G78gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218));
  INV_X1    g017(.A(G71gat), .ZN(new_n219));
  INV_X1    g018(.A(G78gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n217), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n217), .B1(new_n216), .B2(new_n221), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n215), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n224), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT100), .A3(new_n222), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT21), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n214), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n214), .B1(new_n212), .B2(new_n232), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n231), .A2(KEYINPUT21), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI22_X1  g037(.A1(new_n234), .A2(new_n235), .B1(KEYINPUT21), .B2(new_n231), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G231gat), .ZN(new_n241));
  INV_X1    g040(.A(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(new_n242), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G183gat), .B(G211gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT20), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT14), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G29gat), .B2(G36gat), .ZN(new_n256));
  OR3_X1    g055(.A1(new_n255), .A2(G29gat), .A3(G36gat), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT91), .B(G29gat), .Z(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT92), .B(G36gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G43gat), .B(G50gat), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n261), .A2(KEYINPUT15), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n260), .A2(new_n262), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(KEYINPUT15), .B2(new_n261), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT94), .A2(KEYINPUT17), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT94), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT17), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n265), .A2(new_n270), .A3(new_n271), .A4(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G85gat), .A2(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT7), .ZN(new_n277));
  NAND2_X1  g076(.A1(G99gat), .A2(G106gat), .ZN(new_n278));
  INV_X1    g077(.A(G85gat), .ZN(new_n279));
  INV_X1    g078(.A(G92gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(KEYINPUT8), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G99gat), .B(G106gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n283), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n282), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G190gat), .B(G218gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G134gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT102), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n292), .A2(new_n301), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n284), .A2(new_n228), .A3(new_n225), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT10), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n223), .A2(new_n224), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT103), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT103), .A4(new_n308), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(KEYINPUT10), .B(new_n287), .C1(new_n226), .C2(new_n229), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n306), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT104), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n316), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n320), .B1(new_n313), .B2(new_n314), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT104), .B1(new_n321), .B2(new_n306), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n306), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G120gat), .B(G148gat), .Z(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(G204gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT105), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n317), .ZN(new_n333));
  INV_X1    g132(.A(new_n329), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n324), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n254), .A2(new_n304), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT99), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  INV_X1    g139(.A(G64gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(new_n280), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(KEYINPUT23), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n348), .A2(G169gat), .A3(G176gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT24), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(KEYINPUT24), .ZN(new_n353));
  INV_X1    g152(.A(G183gat), .ZN(new_n354));
  INV_X1    g153(.A(G190gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(KEYINPUT23), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n348), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(KEYINPUT64), .A3(new_n359), .A4(new_n345), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n350), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR3_X1   g164(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT23), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n347), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n357), .A2(new_n367), .A3(KEYINPUT25), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n351), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n372), .A2(KEYINPUT67), .A3(new_n345), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT67), .B1(new_n372), .B2(new_n345), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT68), .B(KEYINPUT26), .Z(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n365), .B2(new_n366), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n371), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n355), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(KEYINPUT66), .A3(KEYINPUT28), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT27), .B(G183gat), .ZN(new_n383));
  OR2_X1    g182(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n384));
  NAND2_X1  g183(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n383), .A2(new_n355), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n370), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT75), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n345), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT67), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n372), .A2(KEYINPUT67), .A3(new_n345), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT68), .B(KEYINPUT26), .ZN(new_n398));
  INV_X1    g197(.A(new_n366), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n364), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n351), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT69), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n386), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT69), .B1(new_n378), .B2(new_n387), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n370), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n391), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n363), .A2(new_n369), .B1(new_n378), .B2(new_n387), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n408), .B(new_n390), .C1(new_n409), .C2(KEYINPUT29), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G197gat), .B(G204gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT22), .ZN(new_n413));
  INV_X1    g212(.A(G211gat), .ZN(new_n414));
  INV_X1    g213(.A(G218gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT22), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n412), .B1(new_n420), .B2(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n424), .A3(new_n390), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n391), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n422), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n339), .B(new_n343), .C1(new_n423), .C2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n429), .A3(new_n343), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n423), .A2(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(new_n343), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n339), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(G141gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(G148gat), .ZN(new_n441));
  INV_X1    g240(.A(G148gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(G141gat), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT78), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT2), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT79), .ZN(new_n448));
  INV_X1    g247(.A(G155gat), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n446), .B(new_n448), .C1(new_n449), .C2(new_n295), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n442), .A2(G141gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n440), .A2(G148gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G155gat), .B(G162gat), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G134gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G113gat), .B(G120gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(G127gat), .ZN(new_n463));
  INV_X1    g262(.A(G127gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G134gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI221_X1 g265(.A(new_n461), .B1(new_n462), .B2(KEYINPUT1), .C1(KEYINPUT70), .C2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(G155gat), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT2), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT80), .B1(new_n441), .B2(new_n443), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n451), .A2(new_n452), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n457), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G120gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G113gat), .ZN(new_n477));
  INV_X1    g276(.A(G113gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G120gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT1), .ZN(new_n483));
  XNOR2_X1  g282(.A(G127gat), .B(G134gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT71), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n459), .A2(new_n467), .A3(new_n475), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n483), .A2(new_n480), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n466), .B1(KEYINPUT71), .B2(new_n462), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT1), .B1(new_n480), .B2(new_n481), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n461), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n459), .A4(new_n475), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n459), .A2(new_n475), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT3), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n467), .A2(new_n486), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT3), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n459), .A2(new_n500), .A3(new_n475), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n439), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n439), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n497), .A2(new_n499), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n487), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n497), .A2(KEYINPUT82), .A3(new_n499), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT39), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n503), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G1gat), .B(G29gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT0), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G57gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n279), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n503), .B2(new_n510), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT40), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n496), .A2(new_n439), .A3(new_n502), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n504), .A3(new_n508), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n496), .A2(new_n502), .A3(KEYINPUT5), .A4(new_n439), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n523), .A2(KEYINPUT86), .A3(new_n524), .A4(new_n525), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n516), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n528), .A2(KEYINPUT87), .A3(new_n516), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n511), .A2(new_n517), .A3(KEYINPUT40), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n438), .A2(new_n520), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G22gat), .B(G50gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n421), .A2(KEYINPUT84), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT84), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n412), .B(new_n540), .C1(new_n420), .C2(new_n416), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n539), .A2(new_n419), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n500), .B1(new_n542), .B2(KEYINPUT29), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n497), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n422), .B1(new_n501), .B2(new_n424), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n422), .A2(new_n424), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n549), .A2(new_n500), .B1(new_n459), .B2(new_n475), .ZN(new_n550));
  OAI211_X1 g349(.A(G228gat), .B(G233gat), .C1(new_n545), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n548), .B2(new_n551), .ZN(new_n555));
  XOR2_X1   g354(.A(G78gat), .B(G106gat), .Z(new_n556));
  NOR3_X1   g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(new_n551), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT31), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(new_n553), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n538), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n556), .B1(new_n554), .B2(new_n555), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n553), .A3(new_n558), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n537), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n536), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT6), .B1(new_n526), .B2(new_n515), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n534), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT88), .ZN(new_n571));
  INV_X1    g370(.A(new_n526), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT6), .A3(new_n516), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n534), .A2(new_n574), .A3(new_n569), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n435), .B1(new_n434), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT38), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n425), .A2(new_n422), .A3(new_n426), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n579), .B(KEYINPUT37), .C1(new_n411), .C2(new_n422), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n577), .B1(new_n576), .B2(new_n434), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT38), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n436), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n568), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT76), .B1(new_n430), .B2(new_n432), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n588), .B(new_n431), .C1(new_n436), .C2(new_n339), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n569), .A2(KEYINPUT83), .B1(new_n515), .B2(new_n526), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT83), .ZN(new_n592));
  AOI211_X1 g391(.A(new_n592), .B(KEYINPUT6), .C1(new_n526), .C2(new_n515), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n573), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n594), .A3(new_n437), .ZN(new_n595));
  INV_X1    g394(.A(new_n566), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n406), .A2(new_n493), .ZN(new_n598));
  INV_X1    g397(.A(G227gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n242), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n499), .B(new_n370), .C1(new_n404), .C2(new_n405), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT32), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT73), .ZN(new_n604));
  XNOR2_X1  g403(.A(G15gat), .B(G43gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n219), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G99gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(new_n611), .A3(KEYINPUT32), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n604), .A2(new_n607), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n608), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n602), .A2(KEYINPUT32), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n617));
  INV_X1    g416(.A(new_n600), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT34), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT34), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n613), .A2(new_n623), .A3(new_n615), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT74), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(KEYINPUT74), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n625), .B(new_n626), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n613), .A2(new_n615), .A3(new_n623), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n623), .B1(new_n613), .B2(new_n615), .ZN(new_n632));
  OAI22_X1  g431(.A1(new_n631), .A2(new_n632), .B1(KEYINPUT74), .B2(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n586), .A2(new_n597), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n632), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT89), .B1(new_n636), .B2(new_n566), .ZN(new_n637));
  AND4_X1   g436(.A1(KEYINPUT89), .A2(new_n625), .A3(new_n566), .A4(new_n626), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n590), .A2(new_n594), .A3(KEYINPUT35), .A4(new_n437), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n641));
  INV_X1    g440(.A(new_n636), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n596), .ZN(new_n643));
  INV_X1    g442(.A(new_n438), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT35), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G169gat), .B(G197gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT12), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n275), .A2(new_n209), .ZN(new_n656));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n210), .A2(new_n211), .A3(new_n268), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(KEYINPUT97), .A2(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g459(.A1(KEYINPUT97), .A2(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n655), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n209), .B(new_n665), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n666), .A2(new_n268), .B1(new_n275), .B2(new_n209), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(KEYINPUT18), .A3(new_n657), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n657), .B(KEYINPUT13), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n666), .A2(new_n268), .ZN(new_n671));
  INV_X1    g470(.A(new_n658), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n662), .A2(new_n668), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n664), .B(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n338), .B1(new_n648), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n664), .A2(new_n674), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n664), .A2(new_n674), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(KEYINPUT99), .B(new_n679), .C1(new_n635), .C2(new_n647), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n337), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT106), .B(new_n337), .C1(new_n676), .C2(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n594), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(KEYINPUT16), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n208), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n208), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n685), .A2(new_n438), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g494(.A(new_n644), .B(new_n691), .C1(new_n683), .C2(new_n684), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n685), .A2(new_n438), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n696), .A2(new_n690), .B1(new_n697), .B2(G8gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n698), .B2(new_n694), .ZN(G1325gat));
  AOI21_X1  g498(.A(G15gat), .B1(new_n685), .B2(new_n636), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n634), .B(KEYINPUT107), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n683), .B2(new_n684), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(G15gat), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n596), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT108), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n704), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(new_n258), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n645), .A2(new_n646), .ZN(new_n710));
  INV_X1    g509(.A(new_n640), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n574), .B1(new_n534), .B2(new_n569), .ZN(new_n713));
  INV_X1    g512(.A(new_n569), .ZN(new_n714));
  AOI211_X1 g513(.A(KEYINPUT88), .B(new_n714), .C1(new_n532), .C2(new_n533), .ZN(new_n715));
  INV_X1    g514(.A(new_n573), .ZN(new_n716));
  INV_X1    g515(.A(new_n581), .ZN(new_n717));
  NOR4_X1   g516(.A1(new_n713), .A2(new_n715), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n585), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n567), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n595), .A2(KEYINPUT109), .A3(new_n596), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT109), .B1(new_n595), .B2(new_n596), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n634), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT110), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n634), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n597), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n595), .A2(KEYINPUT109), .A3(new_n596), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n730), .A3(new_n586), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n712), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n304), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n709), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n648), .A2(KEYINPUT44), .A3(new_n304), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n254), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n679), .A3(new_n336), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n708), .B1(new_n739), .B2(new_n594), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n648), .A2(new_n675), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n648), .A2(new_n338), .A3(new_n675), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n733), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n737), .A2(new_n336), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n594), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n741), .B1(new_n748), .B2(new_n258), .ZN(new_n749));
  NOR4_X1   g548(.A1(new_n747), .A2(KEYINPUT45), .A3(new_n594), .A4(new_n708), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(G1328gat));
  NAND4_X1  g550(.A1(new_n745), .A2(new_n259), .A3(new_n438), .A4(new_n746), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n644), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n259), .ZN(G1329gat));
  OAI21_X1  g555(.A(G43gat), .B1(new_n739), .B2(new_n634), .ZN(new_n757));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n745), .A2(new_n758), .A3(new_n636), .A4(new_n746), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(KEYINPUT47), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n701), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n734), .A2(new_n761), .A3(new_n738), .A4(new_n735), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT47), .B1(new_n763), .B2(new_n759), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT111), .B(KEYINPUT47), .C1(new_n763), .C2(new_n759), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(G1330gat));
  NAND4_X1  g567(.A1(new_n734), .A2(new_n596), .A3(new_n738), .A4(new_n735), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G50gat), .ZN(new_n770));
  INV_X1    g569(.A(G50gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n745), .A2(new_n771), .A3(new_n596), .A4(new_n746), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT112), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n773), .B(new_n775), .ZN(G1331gat));
  NOR2_X1   g575(.A1(new_n732), .A2(new_n675), .ZN(new_n777));
  INV_X1    g576(.A(new_n336), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n254), .A2(new_n778), .A3(new_n304), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n686), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g582(.A(new_n438), .B(KEYINPUT114), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n777), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n785), .A2(KEYINPUT115), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1333gat));
  OAI21_X1  g590(.A(new_n219), .B1(new_n780), .B2(new_n642), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n761), .A2(G71gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n780), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n566), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n220), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n737), .A2(new_n675), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n778), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n736), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT116), .B1(new_n801), .B2(new_n594), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n736), .A2(new_n803), .A3(new_n686), .A4(new_n800), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(G85gat), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NOR4_X1   g605(.A1(new_n732), .A2(new_n806), .A3(new_n733), .A4(new_n799), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n724), .A2(new_n731), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n647), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n304), .A3(new_n798), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n806), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n336), .A2(new_n279), .A3(new_n686), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n805), .B1(new_n814), .B2(new_n815), .ZN(G1336gat));
  NAND3_X1  g615(.A1(new_n784), .A2(new_n336), .A3(new_n280), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT117), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n733), .B1(new_n809), .B2(new_n647), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n819), .B2(new_n798), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n807), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n734), .A2(new_n735), .A3(new_n784), .A4(new_n800), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G92gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n734), .A2(new_n438), .A3(new_n735), .A4(new_n800), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G92gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n824), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT118), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n813), .A2(new_n818), .B1(G92gat), .B2(new_n826), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n824), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(G1337gat));
  OAI21_X1  g633(.A(G99gat), .B1(new_n801), .B2(new_n701), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n778), .A2(G99gat), .A3(new_n642), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n814), .B2(new_n836), .ZN(G1338gat));
  NAND3_X1  g636(.A1(new_n736), .A2(new_n596), .A3(new_n800), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n778), .A2(G106gat), .A3(new_n566), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n813), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1339gat));
  OR2_X1    g645(.A1(new_n674), .A2(new_n654), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n667), .A2(new_n657), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n671), .A2(new_n672), .A3(new_n670), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n653), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n336), .ZN(new_n853));
  INV_X1    g652(.A(new_n335), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  INV_X1    g654(.A(new_n322), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n321), .A2(KEYINPUT104), .A3(new_n306), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n321), .A2(new_n306), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n333), .A2(KEYINPUT54), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n329), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n319), .A2(new_n322), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n334), .B1(new_n863), .B2(new_n855), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n854), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n675), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n304), .B1(new_n853), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n864), .B2(new_n860), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n865), .A2(new_n858), .A3(new_n329), .A4(new_n860), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n335), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n733), .A2(new_n872), .A3(new_n851), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n254), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n337), .A2(new_n679), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n643), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n594), .A3(new_n784), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n679), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n594), .B1(new_n874), .B2(new_n875), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n637), .A2(new_n638), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n784), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n478), .A3(new_n675), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n880), .A2(new_n886), .ZN(G1340gat));
  AOI21_X1  g686(.A(new_n476), .B1(new_n878), .B2(new_n336), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT119), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n476), .A3(new_n336), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1341gat));
  AOI21_X1  g690(.A(G127gat), .B1(new_n885), .B2(new_n737), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n254), .A2(new_n464), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n878), .B2(new_n893), .ZN(G1342gat));
  NOR2_X1   g693(.A1(new_n733), .A2(new_n438), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n883), .A2(new_n460), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT56), .Z(new_n897));
  OAI21_X1  g696(.A(G134gat), .B1(new_n879), .B2(new_n733), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n679), .A2(G141gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n701), .A2(new_n596), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT121), .Z(new_n902));
  AND2_X1   g701(.A1(new_n902), .A2(new_n881), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT123), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n902), .A2(KEYINPUT123), .A3(new_n881), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n884), .B(new_n900), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n254), .A2(new_n675), .A3(new_n304), .A4(new_n336), .ZN(new_n907));
  INV_X1    g706(.A(new_n873), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n851), .B1(new_n335), .B2(new_n332), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n679), .B1(new_n872), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n867), .A2(KEYINPUT120), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n913), .B2(new_n304), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n914), .B2(new_n254), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT57), .B1(new_n915), .B2(new_n566), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n566), .B1(new_n874), .B2(new_n875), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n725), .A2(new_n784), .A3(new_n594), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G141gat), .B1(new_n921), .B2(new_n679), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n884), .A3(new_n900), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n903), .A2(KEYINPUT122), .A3(new_n884), .A4(new_n900), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n927), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n929), .B2(new_n923), .ZN(G1344gat));
  NAND2_X1  g729(.A1(new_n902), .A2(new_n881), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT123), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n884), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n336), .A2(new_n442), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(new_n921), .B2(new_n778), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n442), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n918), .B1(new_n915), .B2(new_n566), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n917), .A2(KEYINPUT57), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n336), .A3(new_n920), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n936), .B1(new_n942), .B2(G148gat), .ZN(new_n943));
  OAI22_X1  g742(.A1(new_n934), .A2(new_n935), .B1(new_n938), .B2(new_n943), .ZN(G1345gat));
  NOR3_X1   g743(.A1(new_n921), .A2(new_n449), .A3(new_n254), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n933), .A2(new_n737), .A3(new_n884), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n449), .ZN(G1346gat));
  OAI211_X1 g746(.A(new_n468), .B(new_n469), .C1(new_n921), .C2(new_n733), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n468), .A2(new_n469), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n895), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n932), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n948), .B(new_n953), .C1(new_n932), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n644), .A2(new_n686), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n876), .A2(new_n643), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957), .B2(new_n679), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n884), .B1(new_n874), .B2(new_n875), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n594), .A3(new_n882), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n679), .A2(G169gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1348gat));
  OAI21_X1  g761(.A(G176gat), .B1(new_n957), .B2(new_n778), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n778), .A2(G176gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT125), .Z(G1349gat));
  OAI21_X1  g765(.A(G183gat), .B1(new_n957), .B2(new_n254), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n737), .A2(new_n383), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g769(.A(G190gat), .B1(new_n957), .B2(new_n733), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n304), .A2(new_n355), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n960), .B2(new_n973), .ZN(G1351gat));
  OAI21_X1  g773(.A(new_n675), .B1(new_n867), .B2(KEYINPUT120), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n872), .A2(new_n910), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n853), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n873), .B1(new_n977), .B2(new_n733), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n875), .B1(new_n978), .B2(new_n737), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT57), .B1(new_n979), .B2(new_n596), .ZN(new_n980));
  AOI211_X1 g779(.A(new_n918), .B(new_n566), .C1(new_n874), .C2(new_n875), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n983), .B1(new_n939), .B2(new_n940), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n701), .A2(new_n956), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n985), .A2(new_n986), .A3(new_n675), .A4(new_n987), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT126), .B1(new_n980), .B2(new_n981), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n939), .A2(new_n983), .A3(new_n940), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n675), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n988), .A2(G197gat), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n959), .A2(new_n594), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n994), .A2(new_n901), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  OR3_X1    g795(.A1(new_n996), .A2(G197gat), .A3(new_n679), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n993), .A2(new_n997), .ZN(G1352gat));
  NAND3_X1  g797(.A1(new_n995), .A2(new_n328), .A3(new_n336), .ZN(new_n999));
  XOR2_X1   g798(.A(new_n999), .B(KEYINPUT62), .Z(new_n1000));
  AND3_X1   g799(.A1(new_n985), .A2(new_n336), .A3(new_n987), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n1001), .B2(new_n328), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n995), .A2(new_n414), .A3(new_n737), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n941), .A2(new_n737), .A3(new_n987), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  NAND4_X1  g806(.A1(new_n985), .A2(G218gat), .A3(new_n304), .A4(new_n987), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n415), .B1(new_n996), .B2(new_n733), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1355gat));
endmodule


