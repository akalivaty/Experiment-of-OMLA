

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594;

  XNOR2_X1 U327 ( .A(n396), .B(n395), .ZN(n578) );
  NOR2_X1 U328 ( .A1(n539), .A2(n468), .ZN(n460) );
  XNOR2_X1 U329 ( .A(n391), .B(KEYINPUT48), .ZN(n552) );
  XNOR2_X1 U330 ( .A(n478), .B(n477), .ZN(n527) );
  XOR2_X1 U331 ( .A(n364), .B(n347), .Z(n295) );
  XNOR2_X1 U332 ( .A(n335), .B(G1GAT), .ZN(n336) );
  XNOR2_X1 U333 ( .A(n337), .B(n336), .ZN(n340) );
  INV_X1 U334 ( .A(G183GAT), .ZN(n319) );
  XNOR2_X1 U335 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U336 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U337 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n477) );
  XNOR2_X1 U338 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U339 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U340 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U341 ( .A(n322), .B(n321), .ZN(n449) );
  XNOR2_X1 U342 ( .A(n355), .B(n354), .ZN(n359) );
  XNOR2_X1 U343 ( .A(n452), .B(n451), .ZN(n539) );
  XNOR2_X1 U344 ( .A(n418), .B(n417), .ZN(n551) );
  XNOR2_X1 U345 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U346 ( .A(n481), .B(G43GAT), .ZN(n482) );
  XNOR2_X1 U347 ( .A(n483), .B(n482), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(G92GAT), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT74), .B(KEYINPUT64), .Z(n299) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G85GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(n301), .B(n300), .Z(n308) );
  XOR2_X1 U355 ( .A(G29GAT), .B(G50GAT), .Z(n303) );
  XNOR2_X1 U356 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n338) );
  XOR2_X1 U358 ( .A(G218GAT), .B(G190GAT), .Z(n305) );
  NAND2_X1 U359 ( .A1(G232GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n338), .B(n306), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n316) );
  XOR2_X1 U363 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n310) );
  XNOR2_X1 U364 ( .A(KEYINPUT73), .B(KEYINPUT11), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U366 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n312) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G162GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(n314), .B(n313), .Z(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n486) );
  XOR2_X1 U371 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n318) );
  XNOR2_X1 U372 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n322) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G176GAT), .ZN(n320) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G8GAT), .Z(n342) );
  XOR2_X1 U376 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n327) );
  XOR2_X1 U377 ( .A(G211GAT), .B(KEYINPUT21), .Z(n324) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n429) );
  XNOR2_X1 U380 ( .A(G204GAT), .B(G92GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n325), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U382 ( .A(n429), .B(n347), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U384 ( .A(n342), .B(n328), .Z(n330) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U387 ( .A(n449), .B(n331), .Z(n462) );
  BUF_X1 U388 ( .A(n462), .Z(n530) );
  XNOR2_X1 U389 ( .A(KEYINPUT122), .B(n530), .ZN(n392) );
  INV_X1 U390 ( .A(n486), .ZN(n564) );
  XOR2_X1 U391 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n333) );
  XNOR2_X1 U392 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n346) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G15GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n334), .B(G113GAT), .ZN(n450) );
  XOR2_X1 U396 ( .A(G141GAT), .B(G22GAT), .Z(n422) );
  XOR2_X1 U397 ( .A(n450), .B(n422), .Z(n337) );
  NAND2_X1 U398 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  XOR2_X1 U399 ( .A(n338), .B(KEYINPUT67), .Z(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G197GAT), .Z(n341) );
  XOR2_X1 U402 ( .A(n346), .B(n345), .Z(n555) );
  XOR2_X1 U403 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n364) );
  NAND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n295), .B(n348), .ZN(n349) );
  XOR2_X1 U406 ( .A(G85GAT), .B(G57GAT), .Z(n397) );
  XNOR2_X1 U407 ( .A(n349), .B(n397), .ZN(n355) );
  XOR2_X1 U408 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n351) );
  XNOR2_X1 U409 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U411 ( .A(G176GAT), .B(KEYINPUT72), .Z(n352) );
  XNOR2_X1 U412 ( .A(G99GAT), .B(G71GAT), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n356), .B(G120GAT), .ZN(n447) );
  XNOR2_X1 U414 ( .A(G106GAT), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n357), .B(G148GAT), .ZN(n427) );
  XOR2_X1 U416 ( .A(n447), .B(n427), .Z(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n586) );
  XNOR2_X1 U418 ( .A(KEYINPUT41), .B(n586), .ZN(n512) );
  NAND2_X1 U419 ( .A1(n555), .A2(n512), .ZN(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n381) );
  XOR2_X1 U422 ( .A(G211GAT), .B(G127GAT), .Z(n363) );
  XNOR2_X1 U423 ( .A(G22GAT), .B(G183GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U425 ( .A(n365), .B(n364), .Z(n367) );
  XNOR2_X1 U426 ( .A(G15GAT), .B(G71GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n380) );
  XOR2_X1 U428 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n369) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U431 ( .A(n370), .B(KEYINPUT77), .Z(n378) );
  XOR2_X1 U432 ( .A(G64GAT), .B(G78GAT), .Z(n372) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(G155GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n374) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(G57GAT), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n589) );
  INV_X1 U441 ( .A(n589), .ZN(n562) );
  NOR2_X1 U442 ( .A1(n381), .A2(n562), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n382), .B(KEYINPUT117), .ZN(n383) );
  NOR2_X1 U444 ( .A1(n564), .A2(n383), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n384), .B(KEYINPUT47), .ZN(n390) );
  XOR2_X1 U446 ( .A(n555), .B(KEYINPUT69), .Z(n567) );
  XNOR2_X1 U447 ( .A(KEYINPUT36), .B(n486), .ZN(n592) );
  NOR2_X1 U448 ( .A1(n592), .A2(n589), .ZN(n385) );
  XNOR2_X1 U449 ( .A(KEYINPUT45), .B(n385), .ZN(n386) );
  NAND2_X1 U450 ( .A1(n386), .A2(n586), .ZN(n387) );
  NOR2_X1 U451 ( .A1(n567), .A2(n387), .ZN(n388) );
  XOR2_X1 U452 ( .A(KEYINPUT118), .B(n388), .Z(n389) );
  NAND2_X1 U453 ( .A1(n390), .A2(n389), .ZN(n391) );
  NAND2_X1 U454 ( .A1(n392), .A2(n552), .ZN(n396) );
  INV_X1 U455 ( .A(KEYINPUT54), .ZN(n394) );
  INV_X1 U456 ( .A(KEYINPUT123), .ZN(n393) );
  XOR2_X1 U457 ( .A(n397), .B(KEYINPUT75), .Z(n400) );
  XNOR2_X1 U458 ( .A(G134GAT), .B(G127GAT), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n398), .B(KEYINPUT0), .ZN(n440) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(n440), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n413) );
  XOR2_X1 U462 ( .A(G148GAT), .B(G120GAT), .Z(n402) );
  XNOR2_X1 U463 ( .A(G113GAT), .B(G141GAT), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U465 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n404) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U468 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n408) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(KEYINPUT91), .B(n409), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U475 ( .A(KEYINPUT3), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U476 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(KEYINPUT87), .B(n416), .Z(n430) );
  INV_X1 U479 ( .A(n430), .ZN(n417) );
  INV_X1 U480 ( .A(n551), .ZN(n577) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n420) );
  XNOR2_X1 U482 ( .A(G50GAT), .B(KEYINPUT89), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U484 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n426) );
  XNOR2_X1 U488 ( .A(G204GAT), .B(KEYINPUT88), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n468) );
  AND2_X1 U494 ( .A1(n577), .A2(n468), .ZN(n435) );
  NAND2_X1 U495 ( .A1(n578), .A2(n435), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n436), .B(KEYINPUT124), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n437), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U498 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U499 ( .A(KEYINPUT84), .B(KEYINPUT80), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U501 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U502 ( .A(KEYINPUT79), .B(KEYINPUT82), .Z(n443) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U505 ( .A(KEYINPUT81), .B(n444), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U507 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U509 ( .A1(n453), .A2(n539), .ZN(n575) );
  NOR2_X1 U510 ( .A1(n486), .A2(n575), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n455) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  NAND2_X1 U514 ( .A1(n539), .A2(n530), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n468), .A2(n458), .ZN(n459) );
  XNOR2_X1 U516 ( .A(KEYINPUT25), .B(n459), .ZN(n465) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(n579) );
  XOR2_X1 U519 ( .A(n462), .B(KEYINPUT27), .Z(n469) );
  INV_X1 U520 ( .A(n469), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n579), .A2(n463), .ZN(n554) );
  XNOR2_X1 U522 ( .A(n554), .B(KEYINPUT95), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT96), .ZN(n489) );
  OR2_X1 U525 ( .A1(n551), .A2(n562), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n489), .A2(n467), .ZN(n473) );
  XOR2_X1 U527 ( .A(n468), .B(KEYINPUT28), .Z(n534) );
  NOR2_X1 U528 ( .A1(n469), .A2(n534), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n470), .A2(n551), .ZN(n541) );
  XOR2_X1 U530 ( .A(n539), .B(KEYINPUT85), .Z(n471) );
  NOR2_X1 U531 ( .A1(n541), .A2(n471), .ZN(n491) );
  AND2_X1 U532 ( .A1(n589), .A2(n491), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n475) );
  INV_X1 U534 ( .A(KEYINPUT101), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n592), .A2(n476), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n567), .A2(n586), .ZN(n494) );
  NOR2_X1 U538 ( .A1(n527), .A2(n494), .ZN(n479) );
  XOR2_X1 U539 ( .A(KEYINPUT103), .B(n479), .Z(n480) );
  XNOR2_X1 U540 ( .A(KEYINPUT38), .B(n480), .ZN(n510) );
  NAND2_X1 U541 ( .A1(n539), .A2(n510), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n481) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT97), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT34), .B(n485), .Z(n496) );
  XOR2_X1 U546 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n488) );
  NAND2_X1 U547 ( .A1(n562), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n493) );
  NOR2_X1 U549 ( .A1(n551), .A2(n489), .ZN(n490) );
  OR2_X1 U550 ( .A1(n491), .A2(n490), .ZN(n492) );
  NAND2_X1 U551 ( .A1(n493), .A2(n492), .ZN(n513) );
  NOR2_X1 U552 ( .A1(n494), .A2(n513), .ZN(n501) );
  NAND2_X1 U553 ( .A1(n501), .A2(n551), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n501), .A2(n530), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U558 ( .A1(n501), .A2(n539), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U560 ( .A(G15GAT), .B(n500), .Z(G1326GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n534), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n505) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(n507) );
  NAND2_X1 U567 ( .A1(n510), .A2(n551), .ZN(n506) );
  XOR2_X1 U568 ( .A(n507), .B(n506), .Z(G1328GAT) );
  NAND2_X1 U569 ( .A1(n510), .A2(n530), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U571 ( .A(G36GAT), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n510), .A2(n534), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U574 ( .A(n555), .ZN(n581) );
  INV_X1 U575 ( .A(n512), .ZN(n570) );
  NAND2_X1 U576 ( .A1(n581), .A2(n512), .ZN(n526) );
  NOR2_X1 U577 ( .A1(n526), .A2(n513), .ZN(n514) );
  XNOR2_X1 U578 ( .A(KEYINPUT108), .B(n514), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n523), .A2(n551), .ZN(n517) );
  XOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT109), .Z(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT42), .B(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n523), .A2(n530), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n519), .ZN(G1333GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n521) );
  NAND2_X1 U587 ( .A1(n539), .A2(n523), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U591 ( .A1(n534), .A2(n523), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(n528), .Z(n535) );
  NAND2_X1 U595 ( .A1(n535), .A2(n551), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n535), .A2(n530), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n539), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(KEYINPUT114), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U603 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NAND2_X1 U606 ( .A1(n539), .A2(n552), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n547), .A2(n567), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U611 ( .A1(n547), .A2(n512), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  NAND2_X1 U613 ( .A1(n547), .A2(n562), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U617 ( .A1(n547), .A2(n564), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U619 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n565), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U626 ( .A1(n565), .A2(n512), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .Z(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U634 ( .A(n567), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n568), .A2(n575), .ZN(n569) );
  XOR2_X1 U636 ( .A(G169GAT), .B(n569), .Z(G1348GAT) );
  NOR2_X1 U637 ( .A1(n575), .A2(n570), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT56), .Z(n572) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NOR2_X1 U642 ( .A1(n589), .A2(n575), .ZN(n576) );
  XOR2_X1 U643 ( .A(G183GAT), .B(n576), .Z(G1350GAT) );
  AND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n591) );
  NOR2_X1 U646 ( .A1(n591), .A2(n581), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  NOR2_X1 U651 ( .A1(n591), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n591), .ZN(n590) );
  XOR2_X1 U655 ( .A(G211GAT), .B(n590), .Z(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

