//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G119), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n187), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n191), .A2(new_n193), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n191), .B2(new_n193), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(KEYINPUT0), .B(G128), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT11), .B1(new_n212), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT64), .A2(G131), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT64), .A2(G131), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n217), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n217), .B2(new_n219), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n211), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(G143), .B2(new_n208), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n228), .A2(new_n229), .B1(new_n207), .B2(new_n209), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n203), .A2(G128), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n215), .B2(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT65), .B1(new_n212), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n215), .A3(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n212), .A2(KEYINPUT66), .A3(G137), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n218), .B1(new_n213), .B2(new_n216), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n222), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n233), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n201), .B1(new_n226), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  AND4_X1   g060(.A1(new_n246), .A2(new_n233), .A3(new_n241), .A4(new_n243), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n230), .A2(new_n232), .B1(new_n242), .B2(new_n222), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n248), .B2(new_n241), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n199), .B2(new_n200), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n191), .A2(new_n193), .ZN(new_n253));
  INV_X1    g067(.A(new_n198), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n191), .A2(new_n193), .A3(new_n198), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n226), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n245), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT73), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n244), .A2(KEYINPUT69), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n248), .A2(new_n246), .A3(new_n241), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n226), .A2(new_n252), .A3(new_n257), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n214), .B1(G134), .B2(new_n215), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n212), .A2(KEYINPUT11), .A3(G137), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n219), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G131), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n243), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(new_n211), .B1(new_n248), .B2(new_n241), .ZN(new_n271));
  OAI22_X1  g085(.A1(new_n264), .A2(new_n265), .B1(new_n201), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n226), .A2(new_n244), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n252), .A2(new_n257), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n260), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n279));
  NOR2_X1   g093(.A1(G237), .A2(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G210), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT26), .B(G101), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n201), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n270), .B2(new_n211), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n262), .A3(new_n263), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n275), .B2(new_n287), .ZN(new_n291));
  AOI211_X1 g105(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n226), .C2(new_n244), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n286), .B(new_n289), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n250), .A2(new_n258), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n284), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n278), .A2(new_n285), .B1(KEYINPUT31), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n293), .A2(new_n297), .A3(new_n294), .A4(new_n284), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n264), .A2(new_n265), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT67), .B1(new_n271), .B2(KEYINPUT30), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n275), .A2(new_n290), .A3(new_n287), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n201), .B1(new_n250), .B2(new_n288), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(KEYINPUT72), .A3(new_n297), .A4(new_n284), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n310), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(new_n312), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT76), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n277), .A2(new_n284), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n261), .A2(new_n274), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n306), .B2(new_n284), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n261), .A2(new_n284), .A3(new_n274), .A4(new_n277), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n293), .A2(new_n294), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n285), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT74), .A4(new_n321), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n262), .A2(new_n263), .A3(new_n226), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n250), .A2(new_n258), .B1(new_n328), .B2(new_n276), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT75), .B1(new_n329), .B2(new_n260), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n276), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n294), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT28), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n336));
  AOI21_X1  g150(.A(G902), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n323), .A2(new_n327), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G472), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n309), .A2(new_n340), .A3(new_n315), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n313), .A2(new_n317), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT9), .B(G234), .ZN(new_n343));
  OAI21_X1  g157(.A(G221), .B1(new_n343), .B2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT84), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G140), .ZN(new_n347));
  INV_X1    g161(.A(G227), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G953), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G104), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(new_n352), .B2(G107), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  AOI21_X1  g173(.A(G101), .B1(new_n352), .B2(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n360), .A3(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT85), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n358), .A2(KEYINPUT85), .A3(new_n364), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n362), .B(new_n211), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n223), .A2(new_n225), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT86), .B1(new_n352), .B2(G107), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n355), .A3(G104), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n371), .A3(new_n357), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G101), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n361), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n208), .A2(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n206), .A2(G146), .ZN(new_n376));
  AND4_X1   g190(.A1(new_n227), .A2(new_n375), .A3(new_n376), .A4(G128), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n231), .A2(G128), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n374), .A2(new_n379), .A3(KEYINPUT10), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n353), .A2(new_n356), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n382), .A2(new_n360), .B1(new_n372), .B2(G101), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n383), .B2(new_n233), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n367), .B(new_n368), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT87), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT10), .B1(new_n374), .B2(new_n379), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n381), .A3(new_n233), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n368), .A4(new_n367), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n393), .A2(new_n359), .B1(new_n210), .B2(new_n205), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n358), .A2(new_n364), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n358), .A2(KEYINPUT85), .A3(new_n364), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n387), .A2(new_n388), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n400), .A2(new_n368), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n351), .B1(new_n392), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n351), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n383), .A2(new_n233), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n374), .A2(new_n379), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n368), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n408), .B(KEYINPUT12), .Z(new_n409));
  AOI21_X1  g223(.A(new_n350), .B1(new_n386), .B2(new_n391), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(KEYINPUT88), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n402), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n412), .A2(G469), .A3(G902), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  INV_X1    g228(.A(G902), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n408), .B(KEYINPUT12), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n392), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n418), .A2(new_n350), .B1(new_n410), .B2(new_n401), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n419), .B2(G469), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n346), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G214), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G210), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT8), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n373), .A2(new_n256), .A3(new_n361), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n194), .B1(new_n192), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT90), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n191), .A2(KEYINPUT5), .A3(new_n193), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n431), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n383), .B1(new_n256), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n428), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G125), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n230), .A2(new_n232), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT89), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n205), .A2(G125), .A3(new_n210), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n230), .A2(new_n232), .A3(new_n442), .A4(new_n438), .ZN(new_n443));
  INV_X1    g257(.A(G224), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G953), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT91), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n440), .A2(new_n441), .A3(new_n443), .A4(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n445), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT7), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n451), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n440), .A2(new_n453), .A3(new_n441), .A4(new_n443), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n437), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n437), .A2(new_n452), .A3(KEYINPUT92), .A4(new_n454), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n383), .A2(new_n435), .A3(new_n256), .ZN(new_n459));
  INV_X1    g273(.A(new_n359), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n460), .A2(new_n461), .B1(new_n199), .B2(new_n200), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n366), .A2(new_n365), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n459), .B(new_n427), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n457), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n466));
  INV_X1    g280(.A(new_n427), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n445), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n415), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n426), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n457), .A2(new_n458), .A3(new_n464), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(new_n415), .A3(new_n425), .A4(new_n474), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n424), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n480));
  INV_X1    g294(.A(G237), .ZN(new_n481));
  INV_X1    g295(.A(G953), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G214), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n206), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n280), .A2(G143), .A3(G214), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT18), .A2(G131), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n483), .A2(new_n206), .ZN(new_n488));
  AOI21_X1  g302(.A(G143), .B1(new_n280), .B2(G214), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT18), .B(G131), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G140), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G125), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n438), .A2(G140), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G146), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n493), .A3(new_n208), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n495), .A2(KEYINPUT93), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT93), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n487), .B(new_n490), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT96), .B(G104), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n492), .A2(KEYINPUT16), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT16), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT79), .A4(KEYINPUT16), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(G146), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT80), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n510), .A3(G146), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n208), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n484), .A2(new_n222), .A3(new_n485), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT94), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n517));
  OAI22_X1  g331(.A1(new_n488), .A2(new_n489), .B1(new_n221), .B2(new_n220), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT94), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n484), .A2(new_n519), .A3(new_n222), .A4(new_n485), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n518), .A2(new_n517), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n499), .B(new_n502), .C1(new_n514), .C2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT19), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT19), .B1(new_n492), .B2(new_n493), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n208), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT95), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(new_n208), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n508), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n499), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n502), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n480), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(G146), .B1(new_n506), .B2(new_n507), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(KEYINPUT80), .B2(new_n508), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n511), .A3(new_n522), .A4(new_n521), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n502), .B1(new_n543), .B2(new_n499), .ZN(new_n544));
  INV_X1    g358(.A(new_n524), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n415), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G475), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n536), .A2(new_n480), .A3(new_n537), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT20), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n540), .B(new_n547), .C1(new_n549), .C2(new_n538), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G478), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT99), .B1(new_n229), .B2(G143), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n206), .A3(G128), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n206), .A2(G128), .ZN(new_n558));
  OAI21_X1  g372(.A(G134), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n556), .ZN(new_n560));
  INV_X1    g374(.A(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n212), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT14), .A4(G122), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(G107), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n188), .A2(new_n190), .A3(G122), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT14), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n187), .A2(G122), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n559), .A2(new_n562), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n567), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT98), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n572), .A3(new_n567), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n355), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n565), .A2(new_n572), .A3(new_n567), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n572), .B1(new_n565), .B2(new_n567), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n576), .A2(new_n577), .A3(G107), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n355), .B1(new_n571), .B2(new_n573), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n562), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT13), .B1(new_n554), .B2(new_n556), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n558), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n582), .A2(KEYINPUT100), .B1(KEYINPUT13), .B2(new_n557), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n581), .B2(new_n558), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n212), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n575), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G217), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n343), .A2(new_n588), .A3(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n562), .ZN(new_n592));
  OAI21_X1  g406(.A(G107), .B1(new_n576), .B2(new_n577), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(new_n574), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT100), .B(new_n561), .C1(new_n557), .C2(KEYINPUT13), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n557), .A2(KEYINPUT13), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n585), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G134), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n594), .A2(new_n598), .B1(new_n574), .B2(new_n569), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n589), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n591), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n553), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n598), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n604), .A2(new_n575), .A3(new_n589), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n589), .B1(new_n604), .B2(new_n575), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n415), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT101), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n591), .A2(new_n600), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n602), .A3(new_n415), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n603), .B1(new_n611), .B2(new_n553), .ZN(new_n612));
  OR2_X1    g426(.A1(KEYINPUT102), .A2(G952), .ZN(new_n613));
  NAND2_X1  g427(.A1(KEYINPUT102), .A2(G952), .ZN(new_n614));
  AOI21_X1  g428(.A(G953), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G234), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n481), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT21), .B(G898), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n415), .B(new_n482), .C1(G234), .C2(G237), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n479), .A2(new_n551), .A3(new_n612), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n422), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n588), .B1(G234), .B2(new_n415), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G119), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G128), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(G128), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(KEYINPUT23), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G110), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT78), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR3_X1    g448(.A1(new_n627), .A2(KEYINPUT77), .A3(G128), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT77), .B1(new_n627), .B2(G128), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n628), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT24), .B(G110), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n514), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n631), .A2(G110), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT81), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n508), .A2(new_n496), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT22), .B(G137), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n482), .A2(G221), .A3(G234), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n641), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n640), .A2(new_n514), .B1(new_n646), .B2(new_n647), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n651), .B(KEYINPUT82), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n653), .B(new_n415), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT25), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n641), .A2(new_n648), .ZN(new_n659));
  INV_X1    g473(.A(new_n655), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(KEYINPUT25), .A3(new_n415), .A4(new_n653), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n626), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n626), .A2(new_n415), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n661), .A2(new_n653), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n342), .A2(new_n624), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G101), .ZN(G3));
  INV_X1    g483(.A(G472), .ZN(new_n670));
  AOI21_X1  g484(.A(G902), .B1(new_n296), .B2(new_n308), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n667), .B(new_n311), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n402), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n390), .B1(new_n400), .B2(new_n368), .ZN(new_n675));
  INV_X1    g489(.A(new_n391), .ZN(new_n676));
  OAI211_X1 g490(.A(KEYINPUT88), .B(new_n351), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n417), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n410), .A2(KEYINPUT88), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n414), .A3(new_n415), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n345), .B1(new_n681), .B2(new_n420), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n479), .A2(new_n622), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n601), .A2(G478), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT33), .B1(new_n591), .B2(new_n600), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n599), .B2(new_n589), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT33), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n599), .B2(new_n589), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n587), .A2(KEYINPUT103), .A3(new_n590), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n689), .A3(new_n690), .A4(KEYINPUT104), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n685), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n415), .A2(G478), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n684), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n683), .A2(new_n698), .A3(new_n551), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n673), .A2(new_n682), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT34), .B(G104), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G6));
  NOR2_X1   g516(.A1(new_n672), .A2(new_n422), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n602), .B1(new_n609), .B2(new_n415), .ZN(new_n704));
  AOI211_X1 g518(.A(KEYINPUT101), .B(G902), .C1(new_n591), .C2(new_n600), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n553), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n603), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n551), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n683), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT35), .B(G107), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G9));
  AOI21_X1  g527(.A(new_n670), .B1(new_n309), .B2(new_n415), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n314), .B1(new_n296), .B2(new_n308), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n660), .A2(KEYINPUT36), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n659), .B(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(new_n665), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n663), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n624), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT37), .B(G110), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G12));
  INV_X1    g538(.A(G900), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n618), .B1(new_n725), .B2(new_n620), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n708), .A2(new_n551), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n422), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n479), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n719), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n342), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G128), .ZN(G30));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n734));
  INV_X1    g548(.A(new_n719), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n708), .A2(new_n550), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(new_n424), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n476), .A2(new_n478), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT38), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n295), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n285), .B2(new_n332), .ZN(new_n742));
  OAI21_X1  g556(.A(G472), .B1(new_n742), .B2(G902), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n313), .A2(new_n317), .A3(new_n341), .A4(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n734), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n726), .B(KEYINPUT39), .Z(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n422), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT40), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n313), .A2(new_n317), .A3(new_n341), .A4(new_n743), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n737), .A3(KEYINPUT106), .A4(new_n739), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT40), .B1(new_n422), .B2(new_n747), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n745), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G143), .ZN(G45));
  AOI211_X1 g569(.A(new_n685), .B(new_n696), .C1(new_n693), .C2(new_n694), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n550), .B(new_n727), .C1(new_n756), .C2(new_n684), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n342), .A2(new_n682), .A3(new_n731), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G146), .ZN(G48));
  NAND2_X1  g574(.A1(new_n681), .A2(new_n346), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n680), .A2(new_n415), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n414), .B1(new_n762), .B2(KEYINPUT107), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n680), .A2(new_n764), .A3(new_n415), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n761), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n342), .A2(new_n667), .A3(new_n699), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT41), .B(G113), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G15));
  NAND4_X1  g583(.A1(new_n342), .A2(new_n667), .A3(new_n710), .A4(new_n766), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G116), .ZN(G18));
  OAI21_X1  g585(.A(KEYINPUT107), .B1(new_n412), .B2(G902), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n765), .A3(G469), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n412), .A2(G902), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n345), .B1(new_n774), .B2(new_n414), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n773), .A2(new_n775), .A3(new_n479), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n719), .A2(new_n708), .A3(new_n550), .A4(new_n621), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n342), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G119), .ZN(G21));
  XNOR2_X1  g593(.A(new_n310), .B(KEYINPUT108), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n300), .A2(new_n307), .B1(KEYINPUT31), .B2(new_n295), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n333), .B1(new_n332), .B2(KEYINPUT28), .ZN(new_n782));
  AOI211_X1 g596(.A(KEYINPUT75), .B(new_n260), .C1(new_n294), .C2(new_n331), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n277), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n285), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n780), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n714), .A2(new_n786), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n479), .A2(new_n708), .A3(new_n550), .A4(new_n622), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n667), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n773), .A2(new_n775), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT109), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n479), .A2(new_n708), .A3(new_n550), .A4(new_n622), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n666), .A2(new_n665), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n658), .A2(new_n662), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n626), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n792), .A2(new_n714), .A3(new_n795), .A4(new_n786), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n766), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G122), .ZN(G24));
  NOR3_X1   g614(.A1(new_n714), .A2(new_n786), .A3(new_n719), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n776), .A2(new_n758), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G125), .ZN(G27));
  NOR2_X1   g617(.A1(new_n738), .A2(new_n424), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n682), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n342), .A2(new_n805), .A3(new_n806), .A4(new_n667), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n805), .A2(new_n758), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n313), .A2(new_n339), .A3(new_n316), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(KEYINPUT110), .A3(new_n667), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT110), .B1(new_n809), .B2(new_n667), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n807), .B1(new_n812), .B2(KEYINPUT42), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  INV_X1    g628(.A(new_n728), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n342), .A2(new_n805), .A3(new_n667), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n212), .ZN(G36));
  INV_X1    g631(.A(new_n416), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n418), .A2(new_n350), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n410), .A2(new_n401), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(KEYINPUT111), .A3(G469), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n822), .B2(new_n821), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT111), .B1(new_n823), .B2(G469), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT46), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT46), .B(new_n818), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n681), .A3(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n346), .A2(new_n831), .A3(new_n746), .A4(new_n804), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n551), .B1(new_n756), .B2(new_n684), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT43), .B1(new_n833), .B2(KEYINPUT112), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT113), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n836), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n834), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n714), .A2(new_n715), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n719), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT44), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT44), .A4(new_n842), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n832), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G137), .ZN(G39));
  INV_X1    g662(.A(new_n342), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n849), .A2(new_n795), .A3(new_n758), .A4(new_n804), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n831), .A2(KEYINPUT47), .A3(new_n346), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT47), .B1(new_n831), .B2(new_n346), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  NAND2_X1  g668(.A1(new_n773), .A2(new_n681), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT49), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n667), .A2(new_n346), .A3(new_n423), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n739), .A2(new_n857), .A3(new_n833), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(KEYINPUT49), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n856), .A2(new_n744), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n668), .A2(new_n700), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n668), .A2(new_n700), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n608), .A2(new_n610), .B1(new_n552), .B2(G478), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT115), .B1(new_n866), .B2(new_n603), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n706), .A2(new_n868), .A3(new_n707), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n424), .B(new_n621), .C1(new_n476), .C2(new_n478), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n870), .A2(new_n551), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n703), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n767), .A2(new_n873), .A3(new_n721), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n770), .A2(new_n778), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n865), .A2(new_n799), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n682), .A2(new_n735), .A3(new_n727), .A4(new_n804), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n870), .A2(new_n550), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n342), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n698), .A2(new_n551), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n787), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n816), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n813), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n802), .A2(new_n732), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT116), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n663), .A2(new_n718), .A3(new_n726), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n682), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT117), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n736), .A2(new_n730), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n682), .A2(new_n893), .A3(new_n889), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n751), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(KEYINPUT52), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n802), .A2(new_n732), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n888), .A2(new_n896), .A3(new_n759), .A4(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n759), .A3(new_n802), .A4(new_n732), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n886), .B2(new_n903), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n703), .A2(new_n872), .B1(new_n624), .B2(new_n720), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n905), .A2(new_n767), .A3(new_n770), .A4(new_n778), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n797), .B1(new_n796), .B2(new_n766), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n714), .A2(new_n786), .A3(new_n795), .ZN(new_n908));
  AND4_X1   g722(.A1(new_n797), .A2(new_n766), .A3(new_n908), .A4(new_n788), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(new_n813), .A3(new_n865), .A4(new_n884), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n900), .B(KEYINPUT52), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT53), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n904), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n770), .A2(new_n778), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(new_n799), .A3(new_n767), .A4(new_n905), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n668), .A2(new_n700), .A3(new_n863), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n863), .B1(new_n668), .B2(new_n700), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n812), .A2(KEYINPUT42), .ZN(new_n924));
  INV_X1    g738(.A(new_n807), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n884), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n903), .A2(new_n923), .A3(new_n926), .A4(KEYINPUT53), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n917), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n766), .A2(new_n618), .A3(new_n804), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n931), .A2(new_n744), .A3(new_n667), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n881), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n835), .A2(new_n836), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n908), .A2(new_n618), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n776), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n937), .A3(new_n615), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n934), .A2(new_n931), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n811), .B2(new_n810), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(KEYINPUT48), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(KEYINPUT48), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n934), .A2(new_n804), .A3(new_n935), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT118), .Z(new_n945));
  OR2_X1    g759(.A1(new_n851), .A2(new_n852), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n855), .A2(new_n346), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n756), .A2(new_n550), .A3(new_n684), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n932), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n939), .A2(new_n801), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n790), .A2(new_n739), .A3(new_n423), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n936), .A2(KEYINPUT50), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n936), .A2(new_n954), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n953), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n948), .A2(new_n949), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n949), .B1(new_n948), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n943), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n930), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(G952), .A2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n860), .B1(new_n963), .B2(new_n964), .ZN(G75));
  INV_X1    g779(.A(G210), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n966), .B(new_n415), .C1(new_n917), .C2(new_n927), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n469), .A2(new_n471), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n473), .Z(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n967), .A2(KEYINPUT56), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n917), .A2(new_n927), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(G210), .A3(G902), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT56), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n482), .A2(G952), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n971), .A2(new_n976), .A3(new_n977), .ZN(G51));
  XNOR2_X1  g792(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n416), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n917), .A2(new_n927), .A3(new_n928), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n928), .B1(new_n917), .B2(new_n927), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n680), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n825), .A2(new_n826), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT120), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n973), .A2(G902), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n977), .B1(new_n984), .B2(new_n987), .ZN(G54));
  AND2_X1   g802(.A1(KEYINPUT58), .A2(G475), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n973), .A2(G902), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT121), .ZN(new_n991));
  INV_X1    g805(.A(new_n536), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n990), .B2(new_n992), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n973), .A2(G902), .A3(new_n536), .A4(new_n989), .ZN(new_n995));
  INV_X1    g809(.A(new_n977), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(G60));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n695), .B1(new_n930), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n695), .A2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n981), .B2(new_n982), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n996), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1002), .A2(new_n1005), .ZN(G63));
  NAND2_X1  g820(.A1(G217), .A2(G902), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT60), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n973), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT122), .ZN(new_n1011));
  INV_X1    g825(.A(new_n666), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1008), .B1(new_n917), .B2(new_n927), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT122), .B1(new_n1014), .B2(new_n666), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n977), .B1(new_n1014), .B2(new_n717), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(KEYINPUT61), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT61), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n973), .A2(new_n717), .A3(new_n1009), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n996), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1014), .A2(new_n666), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1017), .A2(new_n1022), .ZN(G66));
  NOR3_X1   g837(.A1(new_n619), .A2(new_n444), .A3(new_n482), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(new_n923), .B2(new_n482), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n968), .B1(G898), .B2(new_n482), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(G69));
  OAI21_X1  g841(.A(G953), .B1(new_n348), .B2(new_n725), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT125), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n849), .A2(new_n795), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n550), .B1(new_n867), .B2(new_n869), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n1031), .A2(new_n881), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1030), .A2(new_n748), .A3(new_n804), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n847), .A2(new_n853), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n888), .A2(new_n759), .A3(new_n898), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n1036), .B2(new_n754), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n759), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n887), .B2(KEYINPUT116), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1040), .A2(new_n754), .A3(new_n1035), .A4(new_n898), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(KEYINPUT124), .ZN(new_n1042));
  AOI21_X1  g856(.A(G953), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n304), .A2(new_n289), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT123), .Z(new_n1045));
  OR2_X1    g859(.A1(new_n525), .A2(new_n526), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1045), .B(new_n1046), .Z(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n831), .A2(new_n346), .A3(new_n746), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n892), .B1(new_n810), .B2(new_n811), .ZN(new_n1051));
  OR2_X1    g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(new_n816), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1036), .A2(new_n1052), .A3(new_n813), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n847), .A2(new_n853), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n482), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n482), .A2(G900), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1047), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1029), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1059), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1029), .ZN(new_n1062));
  OAI211_X1 g876(.A(new_n1061), .B(new_n1062), .C1(new_n1043), .C2(new_n1048), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1060), .A2(new_n1063), .ZN(G72));
  XNOR2_X1  g878(.A(new_n306), .B(KEYINPUT127), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1054), .A2(new_n1055), .A3(new_n877), .ZN(new_n1066));
  XNOR2_X1  g880(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n670), .A2(new_n415), .ZN(new_n1068));
  XOR2_X1   g882(.A(new_n1067), .B(new_n1068), .Z(new_n1069));
  INV_X1    g883(.A(new_n1069), .ZN(new_n1070));
  OAI211_X1 g884(.A(new_n285), .B(new_n1065), .C1(new_n1066), .C2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g885(.A1(new_n904), .A2(new_n915), .ZN(new_n1072));
  INV_X1    g886(.A(new_n326), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1069), .B1(new_n1073), .B2(new_n741), .ZN(new_n1074));
  OAI211_X1 g888(.A(new_n1071), .B(new_n996), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n1038), .A2(new_n1042), .A3(new_n923), .ZN(new_n1076));
  AOI211_X1 g890(.A(new_n285), .B(new_n1065), .C1(new_n1076), .C2(new_n1069), .ZN(new_n1077));
  NOR2_X1   g891(.A1(new_n1075), .A2(new_n1077), .ZN(G57));
endmodule


