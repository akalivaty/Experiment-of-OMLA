//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G113), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n471), .B2(new_n468), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G113), .A3(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n472), .B(new_n474), .C1(new_n466), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  OR2_X1    g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n480), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(G136), .B2(new_n467), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n464), .B2(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n465), .C2(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G114), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n483), .A2(G126), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n496), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n496), .B2(new_n504), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n511), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n509), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n517), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n520), .A2(G89), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n514), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n516), .B1(new_n536), .B2(KEYINPUT73), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n537), .B1(KEYINPUT73), .B2(new_n536), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT74), .B(G90), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n520), .A2(new_n539), .B1(new_n522), .B2(G52), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AND2_X1   g118(.A1(new_n514), .A2(G56), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n520), .A2(G81), .B1(new_n522), .B2(G43), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT77), .Z(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT78), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n534), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(G91), .B2(new_n520), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n522), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  OR2_X1    g141(.A1(new_n517), .A2(new_n524), .ZN(G303));
  NAND2_X1  g142(.A1(new_n520), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n522), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n520), .A2(G86), .B1(new_n522), .B2(G48), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n511), .B2(new_n513), .ZN(new_n574));
  AND2_X1   g149(.A1(G73), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n520), .A2(G85), .B1(new_n522), .B2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n516), .B2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(new_n520), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n534), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(G171), .B2(new_n588), .ZN(G284));
  XOR2_X1   g165(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g166(.A1(G299), .A2(new_n588), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n588), .B2(G168), .ZN(G297));
  OAI21_X1  g168(.A(new_n592), .B1(new_n588), .B2(G168), .ZN(G280));
  INV_X1    g169(.A(new_n587), .ZN(new_n595));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n551), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g177(.A(KEYINPUT3), .B(G2104), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n469), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  INV_X1    g181(.A(G2100), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n467), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n483), .A2(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n480), .A2(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G2096), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n608), .A2(new_n609), .A3(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G2427), .B(G2430), .Z(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(new_n632), .A3(G14), .ZN(G401));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n634));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT17), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(new_n607), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n637), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(new_n615), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(G227));
  XNOR2_X1  g220(.A(G1971), .B(G1976), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT19), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1961), .B(G1966), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n648), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n650), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n657), .C1(new_n647), .C2(new_n656), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G229));
  INV_X1    g239(.A(KEYINPUT24), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G34), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(G34), .ZN(new_n667));
  AOI21_X1  g242(.A(G29), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n478), .B2(G29), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT89), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G2084), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT90), .Z(new_n672));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G33), .ZN(new_n674));
  NAND2_X1  g249(.A1(G115), .A2(G2104), .ZN(new_n675));
  INV_X1    g250(.A(G127), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(new_n466), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n480), .B1(new_n677), .B2(KEYINPUT87), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(KEYINPUT87), .B2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n680));
  NAND2_X1  g255(.A1(G103), .A2(G2104), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(G2105), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n480), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n467), .A2(G139), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n674), .B1(new_n686), .B2(new_n673), .ZN(new_n687));
  OAI21_X1  g262(.A(KEYINPUT94), .B1(G29), .B2(G32), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n467), .A2(G141), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT92), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n469), .A2(G105), .ZN(new_n691));
  NAND3_X1  g266(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT26), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n691), .B(new_n693), .C1(G129), .C2(new_n483), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n690), .A2(KEYINPUT93), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT93), .B1(new_n690), .B2(new_n694), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n695), .A2(new_n696), .A3(new_n673), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n688), .B(KEYINPUT94), .S(new_n697), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT27), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n672), .B1(G2072), .B2(new_n687), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n687), .A2(G2072), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT91), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT96), .ZN(new_n706));
  MUX2_X1   g281(.A(G6), .B(G305), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G23), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT84), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G288), .B2(new_n710), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n709), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n467), .A2(G131), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n483), .A2(G119), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n480), .A2(G107), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G25), .B(new_n727), .S(G29), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(G290), .A2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G24), .ZN(new_n732));
  OR3_X1    g307(.A1(new_n732), .A2(KEYINPUT83), .A3(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT83), .B1(new_n732), .B2(G16), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1986), .Z(new_n736));
  NAND4_X1  g311(.A1(new_n721), .A2(new_n722), .A3(new_n730), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT85), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n673), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n673), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT98), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n710), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n551), .B2(new_n710), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n699), .A2(new_n701), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n670), .A2(G2084), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  NAND4_X1  g328(.A1(new_n747), .A2(new_n750), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n710), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n595), .B2(new_n710), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1348), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n710), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n710), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(G1966), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  OR2_X1    g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  NAND2_X1  g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n762), .A2(new_n673), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n614), .B2(new_n673), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n757), .A2(new_n760), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n467), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n483), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n480), .A2(G116), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n673), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT86), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n673), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n673), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2078), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n710), .A2(G20), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT99), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT23), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n710), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n710), .ZN(new_n791));
  INV_X1    g366(.A(G1961), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n767), .A2(new_n779), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n746), .A2(new_n754), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n706), .A2(new_n740), .A3(new_n795), .ZN(G150));
  INV_X1    g371(.A(G150), .ZN(G311));
  AOI22_X1  g372(.A1(new_n520), .A2(G93), .B1(new_n522), .B2(G55), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n516), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT100), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(new_n550), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n550), .B2(new_n800), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT38), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n595), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n807), .A2(new_n808), .A3(G860), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n801), .A2(G860), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT37), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(new_n811), .ZN(G145));
  NAND2_X1  g387(.A1(new_n483), .A2(G130), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n480), .A2(G118), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G142), .B2(new_n467), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n605), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(new_n727), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n695), .A2(new_n696), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(new_n772), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n772), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n496), .A2(new_n504), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(G2105), .B1(new_n497), .B2(G114), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n503), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n493), .B2(new_n495), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n821), .A2(new_n831), .A3(new_n822), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n685), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n686), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n825), .B2(new_n832), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n819), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(new_n686), .ZN(new_n839));
  INV_X1    g414(.A(new_n819), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n839), .B(new_n840), .C1(new_n833), .C2(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n614), .B(new_n478), .Z(new_n843));
  XNOR2_X1  g418(.A(G162), .B(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(G37), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n838), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT101), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n849), .A2(KEYINPUT40), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT40), .B1(new_n849), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(G395));
  NAND2_X1  g429(.A1(new_n801), .A2(new_n588), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n595), .B1(KEYINPUT102), .B2(G299), .ZN(new_n856));
  AND2_X1   g431(.A1(G299), .A2(KEYINPUT102), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n803), .B(new_n598), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(KEYINPUT41), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(KEYINPUT104), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G305), .ZN(new_n868));
  XNOR2_X1  g443(.A(G290), .B(G288), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(KEYINPUT105), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(KEYINPUT105), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT42), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n866), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n855), .B1(new_n876), .B2(new_n588), .ZN(G295));
  OAI21_X1  g452(.A(new_n855), .B1(new_n876), .B2(new_n588), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n879));
  XNOR2_X1  g454(.A(G301), .B(G286), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n803), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n803), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(KEYINPUT107), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(KEYINPUT107), .B2(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n859), .A3(new_n858), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n860), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n882), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n874), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n865), .A2(KEYINPUT106), .A3(new_n889), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n885), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n884), .A2(new_n888), .B1(new_n862), .B2(new_n889), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n874), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n879), .B1(new_n898), .B2(KEYINPUT43), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n885), .A2(new_n891), .A3(new_n893), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n874), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n902), .A2(new_n903), .A3(new_n897), .A4(new_n894), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n900), .B1(new_n899), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n897), .A3(new_n894), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(KEYINPUT43), .B2(new_n908), .ZN(new_n909));
  OAI22_X1  g484(.A1(new_n905), .A2(new_n906), .B1(new_n909), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g485(.A(KEYINPUT127), .ZN(new_n911));
  INV_X1    g486(.A(G8), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n470), .A2(new_n477), .A3(G40), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n915));
  INV_X1    g490(.A(G1384), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n824), .B2(new_n916), .ZN(new_n917));
  AOI211_X1 g492(.A(KEYINPUT110), .B(G1384), .C1(new_n496), .C2(new_n504), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT50), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G2084), .ZN(new_n922));
  INV_X1    g497(.A(new_n495), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n494), .B1(new_n603), .B2(new_n491), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT71), .B1(new_n925), .B2(new_n830), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n496), .A2(new_n504), .A3(new_n505), .ZN(new_n927));
  AOI21_X1  g502(.A(G1384), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n928), .A2(new_n929), .A3(new_n920), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n916), .B1(new_n506), .B2(new_n507), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT111), .B1(new_n931), .B2(KEYINPUT50), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n921), .B(new_n922), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n917), .B2(new_n918), .ZN(new_n935));
  OAI211_X1 g510(.A(KEYINPUT45), .B(new_n916), .C1(new_n506), .C2(new_n507), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n913), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G1966), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n912), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT113), .B(G8), .ZN(new_n941));
  NOR2_X1   g516(.A1(G168), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT51), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(KEYINPUT51), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n933), .B2(new_n939), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(KEYINPUT120), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT120), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n947), .B(new_n941), .C1(new_n933), .C2(new_n939), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n933), .A2(new_n939), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n942), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n954));
  NOR3_X1   g529(.A1(G166), .A2(new_n954), .A3(new_n912), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(G166), .B2(new_n912), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n920), .B(new_n916), .C1(new_n506), .C2(new_n507), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n913), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT110), .B1(new_n831), .B2(G1384), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n824), .A2(new_n915), .A3(new_n916), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n920), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n961), .A2(new_n964), .A3(G2090), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n824), .A2(new_n916), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n913), .B1(new_n966), .B2(new_n934), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n928), .A2(KEYINPUT109), .A3(KEYINPUT45), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n931), .B2(new_n934), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n965), .B1(new_n972), .B2(new_n713), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n959), .B1(new_n973), .B2(new_n941), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n956), .A2(KEYINPUT112), .A3(new_n957), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT112), .B1(new_n956), .B2(new_n957), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n929), .B1(new_n928), .B2(new_n920), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n931), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n980), .A2(new_n744), .A3(new_n921), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT109), .B1(new_n928), .B2(KEYINPUT45), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n931), .A2(new_n970), .A3(new_n934), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(G1971), .B1(new_n984), .B2(new_n968), .ZN(new_n985));
  OAI211_X1 g560(.A(G8), .B(new_n977), .C1(new_n981), .C2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n962), .A2(new_n913), .A3(new_n963), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n572), .A2(new_n989), .A3(new_n576), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n572), .B2(new_n576), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n992), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n995));
  INV_X1    g570(.A(new_n941), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n987), .A2(new_n993), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G288), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G1976), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(G288), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n987), .A2(new_n996), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n987), .A2(new_n996), .A3(new_n999), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT52), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1004), .A3(KEYINPUT52), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n974), .A2(new_n986), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT123), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n974), .A2(new_n986), .A3(KEYINPUT123), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n980), .A2(new_n921), .ZN(new_n1014));
  INV_X1    g589(.A(G2078), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(new_n968), .C1(new_n969), .C2(new_n971), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n792), .A2(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n962), .A2(new_n963), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n914), .B1(new_n1019), .B2(new_n934), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n1015), .A4(new_n936), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n935), .A2(new_n1015), .A3(new_n913), .A4(new_n936), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT121), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1024), .A3(KEYINPUT53), .ZN(new_n1025));
  AOI21_X1  g600(.A(G301), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1012), .A2(new_n1013), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT125), .B1(new_n953), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1003), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1005), .A2(new_n1004), .A3(KEYINPUT52), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n1006), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n972), .A2(new_n713), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n980), .A2(new_n744), .A3(new_n921), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n912), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n1034), .B2(new_n977), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT123), .B1(new_n1035), .B2(new_n974), .ZN(new_n1036));
  AND4_X1   g611(.A1(KEYINPUT123), .A2(new_n974), .A3(new_n986), .A4(new_n1009), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT125), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1026), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1028), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n950), .B1(new_n949), .B2(new_n952), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT126), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n911), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT126), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1043), .B(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(KEYINPUT127), .A3(new_n1041), .A4(new_n1028), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n997), .A2(new_n1000), .A3(new_n998), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n996), .B(new_n987), .C1(new_n1049), .C2(new_n991), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n986), .B2(new_n1031), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT115), .Z(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n945), .A2(G168), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1010), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n958), .B2(new_n1034), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1035), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n967), .B1(new_n982), .B2(new_n983), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n1062), .B2(new_n1015), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1961), .B1(new_n980), .B2(new_n921), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n966), .A2(new_n934), .ZN(new_n1065));
  AND4_X1   g640(.A1(KEYINPUT53), .A2(new_n968), .A3(new_n1015), .A4(new_n1065), .ZN(new_n1066));
  NOR4_X1   g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(G171), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1026), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT122), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n949), .A2(new_n952), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1012), .B(new_n1013), .C1(new_n1068), .C2(KEYINPUT122), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1014), .A2(new_n792), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1025), .A2(new_n1073), .A3(new_n1074), .A4(G301), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT54), .B(new_n1075), .C1(new_n1076), .C2(G301), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT124), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1079));
  OAI21_X1  g654(.A(G171), .B1(new_n1079), .B2(new_n1066), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(KEYINPUT54), .A4(new_n1075), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1071), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n914), .B1(new_n928), .B2(new_n920), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1956), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1062), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(G299), .B(KEYINPUT57), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n987), .A2(G2067), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1014), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g671(.A(KEYINPUT116), .B(new_n1092), .C1(new_n1014), .C2(new_n1093), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n587), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n787), .B1(new_n961), .B2(new_n964), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1088), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n972), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1090), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1091), .B1(new_n1098), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n595), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT60), .B(new_n587), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1108), .A2(new_n1109), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT117), .B(G1996), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1062), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1062), .A2(KEYINPUT118), .A3(new_n1111), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n987), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1118), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT59), .B1(new_n1118), .B2(new_n551), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1091), .A2(new_n1103), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1103), .A2(KEYINPUT119), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(KEYINPUT61), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1091), .B(new_n1103), .C1(KEYINPUT119), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1105), .B1(new_n1110), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1060), .B1(new_n1084), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1045), .A2(new_n1048), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1065), .A2(new_n914), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n820), .B(G1996), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n772), .B(new_n778), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n727), .B(new_n729), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G290), .B(G1986), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1132), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1131), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1132), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n820), .B2(new_n1134), .ZN(new_n1142));
  OR3_X1    g717(.A1(new_n1141), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT46), .B1(new_n1141), .B2(G1996), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT47), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1141), .A2(G1986), .A3(G290), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT48), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1137), .B2(new_n1132), .ZN(new_n1149));
  INV_X1    g724(.A(new_n729), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n727), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1135), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(G2067), .B2(new_n772), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1146), .B(new_n1149), .C1(new_n1132), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1140), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g730(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1157));
  INV_X1    g731(.A(new_n851), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n850), .B1(new_n845), .B2(new_n847), .ZN(new_n1159));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n1160), .A2(new_n909), .ZN(G308));
  AND2_X1   g735(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n1162));
  OAI221_X1 g736(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .C1(new_n1162), .C2(new_n907), .ZN(G225));
endmodule


