//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT33), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n211), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n208), .A2(new_n210), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n220), .A2(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n216), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(new_n221), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n225), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n206), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n231), .A2(new_n206), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n235), .A2(new_n209), .A3(new_n215), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT70), .Z(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n220), .A2(new_n221), .B1(new_n242), .B2(new_n222), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n214), .A2(KEYINPUT28), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT27), .B1(new_n213), .B2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT27), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G183gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n250), .B(new_n214), .C1(KEYINPUT68), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n246), .A2(KEYINPUT69), .A3(KEYINPUT28), .A4(new_n214), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G127gat), .B(G134gat), .Z(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262));
  INV_X1    g061(.A(G113gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(G120gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(G113gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n264), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G113gat), .B(G120gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n260), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT73), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n205), .B1(new_n259), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n226), .A2(new_n227), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n216), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n280), .A2(new_n206), .B1(new_n237), .B2(new_n234), .ZN(new_n281));
  INV_X1    g080(.A(new_n258), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(new_n273), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n273), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n288), .A2(new_n239), .A3(KEYINPUT74), .A4(new_n258), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n277), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G227gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n204), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n283), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n233), .A2(new_n238), .B1(new_n257), .B2(new_n244), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT74), .B1(new_n296), .B2(new_n288), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n204), .B(new_n293), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n203), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n293), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n277), .A2(new_n301), .A3(new_n283), .A4(new_n289), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT34), .ZN(new_n303));
  XOR2_X1   g102(.A(G15gat), .B(G43gat), .Z(new_n304));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT34), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n302), .B(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT75), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT33), .B1(new_n311), .B2(new_n298), .ZN(new_n312));
  INV_X1    g111(.A(new_n306), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n298), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT32), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n307), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n317), .B1(new_n307), .B2(new_n314), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n296), .A2(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT77), .ZN(new_n323));
  OAI22_X1  g122(.A1(new_n321), .A2(new_n323), .B1(new_n296), .B2(new_n322), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n326));
  AND2_X1   g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n328), .B(new_n330), .Z(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n259), .A2(new_n323), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n328), .B(new_n330), .ZN(new_n334));
  INV_X1    g133(.A(new_n322), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n333), .B(new_n334), .C1(new_n321), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n339), .B1(new_n332), .B2(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n332), .A2(KEYINPUT30), .A3(new_n336), .A4(new_n339), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT79), .B(G148gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G141gat), .ZN(new_n348));
  INV_X1    g147(.A(G141gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G148gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G155gat), .ZN(new_n352));
  INV_X1    g151(.A(G162gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  XOR2_X1   g159(.A(G141gat), .B(G148gat), .Z(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n354), .A2(new_n356), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n334), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369));
  INV_X1    g168(.A(G228gat), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n368), .A2(new_n369), .B1(new_n370), .B2(new_n292), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G22gat), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  OAI221_X1 g172(.A(new_n373), .B1(new_n370), .B2(new_n292), .C1(new_n368), .C2(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT31), .B(G50gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n368), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n365), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT3), .B1(new_n334), .B2(new_n367), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n382), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n376), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n374), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n377), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n377), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR4_X1   g189(.A1(new_n319), .A2(new_n320), .A3(new_n346), .A4(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n392));
  XOR2_X1   g191(.A(G1gat), .B(G29gat), .Z(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n288), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n363), .A2(new_n364), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n357), .B1(new_n350), .B2(new_n348), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n366), .A3(new_n284), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n379), .B2(new_n284), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n398), .A2(new_n399), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n379), .B(new_n284), .ZN(new_n408));
  INV_X1    g207(.A(new_n399), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n403), .A2(new_n407), .A3(new_n399), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n379), .A2(new_n284), .A3(new_n404), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n380), .B1(new_n274), .B2(new_n275), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n404), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n397), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n392), .B1(new_n417), .B2(KEYINPUT6), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n406), .A2(new_n410), .B1(new_n415), .B2(new_n412), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NOR4_X1   g219(.A1(new_n419), .A2(KEYINPUT83), .A3(new_n420), .A4(new_n397), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n411), .A2(new_n397), .A3(new_n416), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(new_n423), .B2(KEYINPUT81), .ZN(new_n424));
  INV_X1    g223(.A(new_n397), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n379), .A2(new_n284), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n359), .A2(new_n365), .B1(new_n271), .B2(new_n273), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT5), .B1(new_n428), .B2(new_n399), .ZN(new_n429));
  INV_X1    g228(.A(new_n405), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n379), .B1(new_n286), .B2(new_n287), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(KEYINPUT4), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n403), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n409), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n416), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n425), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n438), .A3(new_n397), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n422), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n307), .A2(new_n314), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n316), .ZN(new_n444));
  INV_X1    g243(.A(new_n390), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT82), .B1(new_n419), .B2(new_n397), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(new_n425), .C1(new_n435), .C2(new_n436), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n424), .A2(new_n439), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n346), .B1(new_n449), .B2(new_n422), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n444), .A2(new_n318), .A3(new_n445), .A4(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n391), .A2(new_n442), .B1(KEYINPUT35), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n332), .A2(new_n336), .A3(new_n339), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n418), .A2(new_n421), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n339), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n332), .A2(new_n336), .ZN(new_n457));
  INV_X1    g256(.A(new_n339), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n455), .B1(new_n332), .B2(new_n336), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT38), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n455), .B1(new_n324), .B2(new_n334), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n333), .B1(new_n321), .B2(new_n335), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n334), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT38), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n464), .B(new_n465), .C1(new_n343), .C2(new_n456), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n454), .A2(new_n461), .A3(new_n466), .A4(new_n440), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n399), .B1(new_n415), .B2(new_n403), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT39), .B1(new_n408), .B2(new_n409), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n471));
  INV_X1    g270(.A(new_n413), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n431), .B2(KEYINPUT4), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n409), .B(new_n471), .C1(new_n473), .C2(new_n433), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n470), .A2(KEYINPUT40), .A3(new_n397), .A4(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n397), .C1(new_n468), .C2(new_n469), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n475), .A2(new_n478), .A3(new_n437), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n390), .B1(new_n479), .B2(new_n346), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n467), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n423), .A2(KEYINPUT81), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n420), .A3(new_n439), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n446), .A2(new_n448), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT83), .B1(new_n437), .B2(new_n420), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n417), .A2(new_n392), .A3(KEYINPUT6), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n482), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n390), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n318), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n319), .B2(new_n320), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n202), .B1(new_n452), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n467), .A2(new_n480), .B1(new_n490), .B2(new_n390), .ZN(new_n498));
  INV_X1    g297(.A(new_n493), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT36), .B1(new_n444), .B2(new_n318), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n444), .A2(new_n318), .A3(new_n445), .A4(new_n482), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n502), .A2(KEYINPUT35), .A3(new_n441), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n501), .B(KEYINPUT86), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G29gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(KEYINPUT14), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(KEYINPUT14), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n513), .B(G36gat), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT15), .B(new_n508), .C1(new_n517), .C2(new_n507), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT16), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n522), .A2(G1gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G8gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n527), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n534), .B(KEYINPUT13), .Z(new_n538));
  AND2_X1   g337(.A1(new_n532), .A2(new_n519), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n532), .A2(new_n519), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n530), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n534), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G197gat), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT11), .B(G169gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT12), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n537), .A2(new_n541), .A3(new_n542), .A4(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n541), .A2(new_n549), .A3(new_n542), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n541), .B2(new_n542), .ZN(new_n551));
  INV_X1    g350(.A(new_n537), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n547), .B(KEYINPUT87), .Z(new_n554));
  OAI21_X1  g353(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n497), .A2(new_n505), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n561), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n562), .A2(new_n570), .A3(KEYINPUT89), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT89), .B1(new_n562), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G127gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT89), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n568), .B1(new_n569), .B2(new_n567), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n562), .A2(new_n570), .A3(KEYINPUT89), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n532), .B1(new_n586), .B2(KEYINPUT21), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(new_n352), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n589), .B(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n580), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n580), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT94), .B1(new_n599), .B2(KEYINPUT7), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n603), .A2(new_n604), .A3(G85gat), .A4(G92gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n606), .A3(KEYINPUT7), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n601), .A2(new_n602), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n609), .B1(new_n608), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n521), .A2(new_n529), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n608), .A2(new_n613), .ZN(new_n618));
  INV_X1    g417(.A(new_n609), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n519), .ZN(new_n623));
  NAND3_X1  g422(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n598), .B1(new_n617), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G134gat), .B(G162gat), .Z(new_n627));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n617), .A2(new_n625), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n596), .B(new_n597), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n626), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n620), .A2(new_n585), .A3(new_n584), .A4(new_n621), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n618), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n562), .A2(new_n570), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n608), .A2(new_n613), .A3(new_n644), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n586), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n641), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G120gat), .B(G148gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n647), .B1(new_n618), .B2(new_n645), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n616), .A2(new_n573), .B1(new_n658), .B2(new_n649), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n659), .B2(new_n640), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n640), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT10), .B1(new_n571), .B2(new_n572), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n616), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n659), .B2(new_n643), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT99), .B1(new_n666), .B2(new_n641), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n663), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n662), .B1(new_n670), .B2(new_n657), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n595), .A2(new_n639), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n556), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n486), .A2(new_n489), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n523), .ZN(G1324gat));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND4_X1  g477(.A1(new_n556), .A2(new_n346), .A3(new_n672), .A4(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n673), .B2(new_n482), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT100), .Z(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n319), .A2(new_n320), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n673), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT101), .Z(new_n690));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n499), .B2(new_n500), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n495), .A2(KEYINPUT102), .A3(new_n493), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n673), .A2(new_n686), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n690), .A2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n673), .A2(new_n445), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  XNOR2_X1  g499(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n701));
  INV_X1    g500(.A(new_n663), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n651), .A2(new_n652), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n668), .B1(new_n703), .B2(new_n640), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT99), .B(new_n641), .C1(new_n651), .C2(new_n652), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n657), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n661), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n556), .A2(new_n595), .A3(new_n639), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n674), .A2(new_n506), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n701), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n709), .A2(new_n701), .A3(new_n710), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n693), .A3(new_n498), .ZN(new_n713));
  INV_X1    g512(.A(new_n452), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT105), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n638), .A2(KEYINPUT44), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n497), .A2(new_n505), .A3(new_n639), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n721), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT104), .B1(new_n721), .B2(KEYINPUT44), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n593), .A2(new_n594), .ZN(new_n725));
  INV_X1    g524(.A(new_n555), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n726), .A3(new_n671), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n674), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n711), .B(new_n712), .C1(new_n729), .C2(new_n506), .ZN(G1328gat));
  NAND2_X1  g529(.A1(new_n346), .A2(new_n514), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT46), .B1(new_n709), .B2(new_n731), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n709), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n728), .A2(new_n346), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n514), .ZN(G1329gat));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n728), .A2(new_n694), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n709), .A2(G43gat), .A3(new_n688), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n694), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(G43gat), .A3(new_n743), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n739), .A2(new_n736), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n744), .B2(new_n745), .ZN(G1330gat));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n724), .A2(new_n390), .A3(new_n727), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G50gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(KEYINPUT107), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n709), .A2(G50gat), .A3(new_n445), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n748), .B2(G50gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n750), .B(new_n752), .ZN(G1331gat));
  NOR4_X1   g552(.A1(new_n595), .A2(new_n555), .A3(new_n639), .A4(new_n708), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n717), .A2(new_n718), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n675), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n563), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n482), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT49), .B(G64gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n758), .B2(new_n761), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n755), .B2(new_n695), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n688), .A2(G71gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n755), .A2(new_n445), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g568(.A1(new_n595), .A2(new_n726), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n638), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n715), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n671), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n611), .A3(new_n674), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n770), .A2(new_n708), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT104), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n721), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n784), .B2(new_n720), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n674), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n786), .B2(new_n611), .ZN(G1336gat));
  AOI21_X1  g586(.A(new_n612), .B1(new_n785), .B2(new_n346), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n346), .A2(new_n612), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n775), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT52), .B1(new_n790), .B2(KEYINPUT109), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n724), .A2(new_n346), .A3(new_n778), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796));
  INV_X1    g595(.A(new_n790), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n791), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(new_n800));
  AOI211_X1 g599(.A(KEYINPUT110), .B(new_n790), .C1(new_n794), .C2(G92gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n792), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n799), .A2(new_n802), .ZN(G1337gat));
  AOI21_X1  g602(.A(G99gat), .B1(new_n776), .B2(new_n687), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n694), .A2(G99gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n785), .B2(new_n805), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n785), .A2(G106gat), .A3(new_n390), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n774), .A2(new_n445), .A3(new_n775), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(G106gat), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n809), .B(KEYINPUT53), .Z(G1339gat));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n667), .A2(new_n811), .A3(new_n669), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n703), .B2(new_n640), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n651), .A2(new_n641), .A3(new_n652), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n657), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n812), .A2(new_n815), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n812), .B2(new_n815), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n661), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n555), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n539), .A2(new_n540), .A3(new_n538), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n534), .B1(new_n530), .B2(new_n533), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n546), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n548), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT112), .B1(new_n671), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n708), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n639), .B1(new_n823), .B2(new_n832), .ZN(new_n833));
  AND4_X1   g632(.A1(new_n639), .A2(new_n820), .A3(new_n822), .A4(new_n828), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n595), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n725), .A2(new_n726), .A3(new_n638), .A4(new_n708), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(KEYINPUT113), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n675), .A3(new_n502), .ZN(new_n842));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n555), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n835), .A2(KEYINPUT113), .A3(new_n836), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n835), .B2(new_n836), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n445), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT114), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n674), .A2(new_n848), .A3(new_n687), .A4(new_n482), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n726), .A2(new_n263), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  AOI21_X1  g650(.A(G120gat), .B1(new_n842), .B2(new_n671), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n708), .A2(new_n266), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n849), .B2(new_n853), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n842), .A2(new_n855), .A3(new_n725), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n849), .A2(new_n725), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n855), .ZN(G1342gat));
  INV_X1    g657(.A(G134gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n859), .A3(new_n639), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT56), .Z(new_n861));
  AND2_X1   g660(.A1(new_n849), .A2(new_n639), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n859), .ZN(G1343gat));
  NOR3_X1   g662(.A1(new_n844), .A2(new_n845), .A3(new_n445), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT115), .B1(new_n864), .B2(KEYINPUT57), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n866), .B(new_n867), .C1(new_n841), .C2(new_n445), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n671), .A2(new_n828), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n639), .B1(new_n823), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n595), .B1(new_n870), .B2(new_n834), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n445), .B1(new_n871), .B2(new_n836), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT57), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n865), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n694), .A2(new_n675), .A3(new_n346), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n555), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n874), .A2(new_n878), .A3(new_n555), .A4(new_n875), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(G141gat), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n846), .A2(new_n695), .A3(new_n674), .A4(new_n390), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n726), .A2(G141gat), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT116), .Z(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n884), .A2(new_n482), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n881), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n876), .A2(G141gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n882), .A2(new_n346), .A3(new_n886), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(KEYINPUT58), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n876), .B2(G141gat), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(KEYINPUT117), .A3(new_n881), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n890), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n901), .B(new_n890), .C1(new_n896), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  AND2_X1   g702(.A1(new_n874), .A2(new_n875), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n347), .C1(new_n904), .C2(new_n671), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n864), .A2(new_n867), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n867), .B2(new_n872), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n671), .A3(new_n875), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n482), .A3(new_n888), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n671), .A2(new_n347), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n905), .A2(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1345gat));
  OR2_X1    g712(.A1(new_n911), .A2(new_n595), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n595), .A2(new_n352), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT121), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n914), .A2(new_n352), .B1(new_n904), .B2(new_n916), .ZN(G1346gat));
  OR2_X1    g716(.A1(new_n911), .A2(new_n638), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n638), .A2(new_n353), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n918), .A2(new_n353), .B1(new_n904), .B2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n674), .A2(new_n482), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n688), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n848), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n218), .A3(new_n726), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n841), .A2(new_n674), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n926), .A2(new_n687), .A3(new_n346), .A4(new_n445), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT122), .Z(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n555), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n925), .B1(new_n929), .B2(new_n218), .ZN(G1348gat));
  NOR3_X1   g729(.A1(new_n924), .A2(new_n219), .A3(new_n708), .ZN(new_n931));
  AOI21_X1  g730(.A(G176gat), .B1(new_n928), .B2(new_n671), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT123), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(KEYINPUT123), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1349gat));
  NOR3_X1   g734(.A1(new_n927), .A2(new_n247), .A3(new_n595), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n938), .B1(new_n924), .B2(new_n595), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G183gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n938), .A3(new_n595), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n924), .B2(new_n638), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n214), .A3(new_n639), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  NAND4_X1  g746(.A1(new_n926), .A2(new_n346), .A3(new_n390), .A4(new_n695), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n555), .ZN(new_n950));
  INV_X1    g749(.A(new_n908), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n694), .A2(new_n922), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT126), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n555), .A2(G197gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  NAND2_X1  g755(.A1(new_n908), .A2(new_n671), .ZN(new_n957));
  OAI21_X1  g756(.A(G204gat), .B1(new_n957), .B2(new_n953), .ZN(new_n958));
  OR3_X1    g757(.A1(new_n948), .A2(G204gat), .A3(new_n708), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT127), .B1(new_n959), .B2(KEYINPUT62), .ZN(new_n961));
  OAI221_X1 g760(.A(new_n958), .B1(KEYINPUT62), .B2(new_n959), .C1(new_n960), .C2(new_n961), .ZN(G1353gat));
  OR3_X1    g761(.A1(new_n948), .A2(G211gat), .A3(new_n595), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n908), .A2(new_n725), .A3(new_n952), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n949), .B2(new_n639), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n639), .A2(G218gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n954), .B2(new_n969), .ZN(G1355gat));
endmodule


