//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  OR2_X1    g010(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n207), .B(new_n210), .C1(new_n214), .C2(KEYINPUT22), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(KEYINPUT75), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n208), .A2(new_n209), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n220));
  OAI21_X1  g019(.A(G218gat), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n217), .B1(new_n223), .B2(new_n207), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT85), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n223), .A2(new_n207), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n215), .A2(KEYINPUT75), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n217), .A3(new_n207), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n225), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n206), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n237), .A2(new_n238), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(G141gat), .B(G148gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(G155gat), .B2(G162gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n236), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G155gat), .ZN(new_n246));
  INV_X1    g045(.A(G162gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT2), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT79), .B1(new_n246), .B2(new_n247), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n245), .B(new_n248), .C1(new_n235), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT86), .B1(new_n234), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n229), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n226), .B1(new_n255), .B2(KEYINPUT85), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT29), .B1(new_n256), .B2(new_n231), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n254), .B(new_n251), .C1(new_n257), .C2(new_n206), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n252), .A2(new_n205), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n233), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(G228gat), .B2(G233gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT3), .B1(new_n260), .B2(new_n233), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT80), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n250), .A3(KEYINPUT80), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(G228gat), .B(G233gat), .C1(new_n270), .C2(new_n262), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT31), .B(G50gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n264), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n264), .B2(new_n271), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n204), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n264), .A2(new_n271), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n272), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n264), .A2(new_n271), .A3(new_n273), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n203), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n282));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT82), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G113gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(G113gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(KEYINPUT71), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(KEYINPUT71), .B2(new_n288), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G127gat), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT1), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n291), .B2(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n293), .B2(G127gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n291), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G120gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n288), .B2(new_n305), .ZN(new_n310));
  OAI211_X1 g109(.A(KEYINPUT70), .B(new_n303), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n304), .A2(G120gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT69), .B1(new_n313), .B2(new_n287), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(new_n308), .A3(new_n307), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT70), .B1(new_n315), .B2(new_n303), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n252), .B(new_n296), .C1(new_n312), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n296), .B1(new_n312), .B2(new_n316), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n267), .A2(KEYINPUT3), .A3(new_n268), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n261), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n311), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n326), .A2(KEYINPUT4), .A3(new_n252), .A4(new_n296), .ZN(new_n327));
  AND4_X1   g126(.A1(new_n285), .A2(new_n319), .A3(new_n322), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n325), .A2(new_n311), .B1(new_n290), .B2(new_n295), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n317), .B1(new_n330), .B2(new_n269), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n284), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n319), .A2(new_n322), .A3(new_n285), .A4(new_n327), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n329), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n282), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G1gat), .B(G29gat), .Z(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n319), .A2(new_n327), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(KEYINPUT5), .A3(new_n285), .A4(new_n322), .ZN(new_n344));
  INV_X1    g143(.A(new_n268), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT80), .B1(new_n242), .B2(new_n250), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n320), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n285), .B1(new_n348), .B2(new_n317), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n334), .B1(new_n329), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n350), .A3(KEYINPUT87), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n342), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n350), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT6), .B1(new_n353), .B2(new_n341), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT66), .B(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n357), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n356), .A2(new_n357), .B1(G190gat), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT23), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n366), .A2(new_n369), .A3(new_n368), .ZN(new_n373));
  INV_X1    g172(.A(new_n361), .ZN(new_n374));
  NAND3_X1  g173(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n374), .B(new_n375), .C1(G183gat), .C2(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT27), .B(G183gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n356), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT28), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n380), .A3(KEYINPUT28), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n365), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT26), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n369), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n365), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n379), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n392), .ZN(new_n394));
  INV_X1    g193(.A(new_n384), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT28), .B1(new_n356), .B2(new_n380), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT25), .B1(new_n373), .B2(new_n376), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n370), .B1(new_n360), .B2(new_n363), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n394), .B1(new_n400), .B2(new_n233), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n259), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n392), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n394), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n260), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT37), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT88), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n402), .A2(new_n405), .A3(new_n409), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n393), .A2(new_n401), .A3(new_n259), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n260), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT76), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT37), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT77), .ZN(new_n419));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n411), .A2(new_n417), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT38), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n344), .A2(new_n350), .A3(KEYINPUT6), .A4(new_n342), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n402), .A2(new_n405), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n422), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n421), .B(KEYINPUT78), .Z(new_n428));
  INV_X1    g227(.A(KEYINPUT38), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n411), .B2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n355), .A2(new_n424), .A3(new_n425), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n343), .A2(new_n322), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n284), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n348), .A2(new_n285), .A3(new_n317), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT39), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT39), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n438), .A3(new_n284), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n341), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT30), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n415), .A2(new_n416), .A3(new_n428), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n426), .B2(new_n422), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n437), .A2(KEYINPUT40), .A3(new_n341), .A4(new_n439), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n447), .A3(new_n352), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n281), .A2(new_n433), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n344), .A2(new_n350), .A3(new_n342), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n344), .A2(new_n350), .A3(KEYINPUT84), .A4(new_n342), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n354), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n425), .ZN(new_n456));
  INV_X1    g255(.A(new_n447), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n276), .A2(new_n280), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n330), .A2(new_n400), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n320), .A2(new_n391), .ZN(new_n462));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n463), .B(KEYINPUT64), .Z(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n472), .A2(KEYINPUT72), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(KEYINPUT72), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT33), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(KEYINPUT32), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n462), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n463), .ZN(new_n481));
  AOI211_X1 g280(.A(KEYINPUT34), .B(new_n464), .C1(new_n461), .C2(new_n462), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n473), .A3(new_n477), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n478), .A2(new_n483), .A3(KEYINPUT73), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n492), .B2(KEYINPUT36), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n450), .A2(new_n460), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n276), .A2(new_n280), .A3(new_n487), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT35), .B1(new_n458), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n443), .A2(new_n444), .A3(new_n497), .A4(new_n446), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n355), .B2(new_n425), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n281), .A2(new_n499), .A3(new_n492), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n494), .B2(new_n501), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(G1gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(G1gat), .B2(new_n506), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G8gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  AOI21_X1  g314(.A(G36gat), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n512), .A2(new_n517), .A3(G29gat), .ZN(new_n518));
  OR3_X1    g317(.A1(new_n516), .A2(KEYINPUT15), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT15), .B1(new_n516), .B2(new_n518), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n520), .B2(new_n521), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n511), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n510), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n505), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n526), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n527), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n523), .B(new_n510), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n529), .B(KEYINPUT13), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G113gat), .B(G141gat), .Z(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT90), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT11), .B(G169gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT12), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n536), .B(new_n542), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n503), .A2(new_n504), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n456), .ZN(new_n545));
  XOR2_X1   g344(.A(G57gat), .B(G64gat), .Z(new_n546));
  NAND2_X1  g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n547), .A2(new_n552), .B1(new_n549), .B2(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n547), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(new_n551), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n546), .B(new_n549), .C1(new_n556), .C2(KEYINPUT91), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n510), .B1(new_n560), .B2(KEYINPUT21), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT93), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G155gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n562), .B(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n558), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(new_n291), .ZN(new_n569));
  XOR2_X1   g368(.A(G183gat), .B(G211gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT41), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT94), .Z(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n576), .A2(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT95), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT96), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n586), .A2(new_n595), .A3(new_n591), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(KEYINPUT97), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n586), .A2(new_n598), .A3(new_n595), .A4(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n583), .B1(new_n600), .B2(new_n523), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n599), .B(new_n597), .C1(new_n524), .C2(new_n525), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n582), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n607), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n581), .A3(new_n605), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n575), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n594), .A2(new_n558), .A3(new_n596), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n614), .B(new_n615), .C1(new_n600), .C2(new_n558), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G230gat), .ZN(new_n619));
  INV_X1    g418(.A(G233gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n615), .B1(new_n600), .B2(new_n558), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n621), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n623), .B2(new_n625), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n613), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n544), .A2(new_n545), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g435(.A1(new_n544), .A2(new_n634), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n637), .A2(KEYINPUT98), .A3(new_n457), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT98), .B1(new_n637), .B2(new_n457), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(G8gat), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n637), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(KEYINPUT42), .A3(new_n447), .A4(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n638), .B2(new_n639), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n640), .B(new_n643), .C1(new_n645), .C2(KEYINPUT42), .ZN(G1325gat));
  AOI21_X1  g445(.A(G15gat), .B1(new_n641), .B2(new_n492), .ZN(new_n647));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n493), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT99), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n641), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n637), .A2(new_n281), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n575), .A2(new_n612), .A3(new_n633), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n544), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n545), .A2(new_n513), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n657), .A2(new_n655), .A3(new_n658), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n447), .B1(new_n455), .B2(new_n425), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n281), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n458), .A2(KEYINPUT101), .A3(new_n459), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n450), .A3(new_n665), .A4(new_n493), .ZN(new_n666));
  AOI211_X1 g465(.A(new_n612), .B(new_n661), .C1(new_n666), .C2(new_n501), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n494), .A2(new_n501), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT89), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n611), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n667), .B1(new_n671), .B2(KEYINPUT44), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n574), .B(KEYINPUT100), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n542), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n536), .B(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n676), .A3(new_n632), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n672), .A2(new_n456), .A3(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n678), .B2(KEYINPUT103), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n659), .B(new_n660), .C1(new_n679), .C2(new_n680), .ZN(G1328gat));
  NAND2_X1  g480(.A1(new_n447), .A2(new_n517), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n657), .A2(KEYINPUT46), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT46), .B1(new_n657), .B2(new_n682), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n672), .A2(new_n457), .A3(new_n677), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n683), .B(new_n684), .C1(new_n685), .C2(new_n517), .ZN(G1329gat));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n672), .A2(new_n493), .A3(new_n677), .ZN(new_n688));
  INV_X1    g487(.A(G43gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  INV_X1    g492(.A(new_n492), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n657), .A2(G43gat), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n690), .B(new_n691), .C1(new_n693), .C2(new_n695), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1330gat));
  INV_X1    g498(.A(G50gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n672), .A2(new_n677), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n459), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n657), .A2(G50gat), .A3(new_n281), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1331gat));
  NAND2_X1  g506(.A1(new_n666), .A2(new_n501), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n613), .A2(new_n676), .A3(new_n632), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n708), .A2(KEYINPUT105), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n456), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g515(.A1(new_n714), .A2(new_n457), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(G1333gat));
  INV_X1    g520(.A(G71gat), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n714), .A2(new_n722), .A3(new_n493), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n712), .A2(new_n492), .A3(new_n713), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  AOI21_X1  g524(.A(G71gat), .B1(new_n724), .B2(KEYINPUT106), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n727), .B(new_n728), .Z(G1334gat));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n281), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g530(.A1(new_n575), .A2(new_n676), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n633), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n672), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n456), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n612), .B1(new_n666), .B2(new_n501), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n732), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n732), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n737), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n741), .A2(KEYINPUT108), .A3(new_n743), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n633), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n545), .A2(new_n588), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n736), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n633), .A2(new_n589), .A3(new_n447), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT110), .Z(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n741), .B2(new_n743), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n589), .B1(new_n734), .B2(new_n447), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n755), .A2(new_n756), .A3(new_n752), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n752), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n735), .B2(new_n493), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n694), .A2(G99gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n747), .B2(new_n761), .ZN(G1338gat));
  INV_X1    g561(.A(new_n733), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n503), .A2(new_n504), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n611), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n459), .B(new_n763), .C1(new_n766), .C2(new_n667), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G106gat), .ZN(new_n768));
  INV_X1    g567(.A(G106gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n633), .A2(new_n769), .A3(new_n459), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n741), .B2(new_n743), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT53), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n768), .B(new_n773), .C1(new_n772), .C2(new_n771), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n770), .B(KEYINPUT111), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n742), .B2(new_n744), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n775), .B(new_n776), .C1(new_n768), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n672), .A2(new_n281), .A3(new_n733), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n769), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n782), .B2(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n774), .B1(new_n780), .B2(new_n783), .ZN(G1339gat));
  NOR3_X1   g583(.A1(new_n613), .A2(new_n676), .A3(new_n633), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n541), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n533), .A2(new_n534), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n529), .B1(new_n526), .B2(new_n527), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(KEYINPUT115), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n787), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n536), .A2(new_n675), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n616), .A2(new_n621), .A3(new_n617), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n621), .B1(new_n616), .B2(new_n617), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  AOI211_X1 g600(.A(KEYINPUT54), .B(new_n621), .C1(new_n616), .C2(new_n617), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n628), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n618), .A2(new_n799), .A3(new_n622), .ZN(new_n804));
  INV_X1    g603(.A(new_n628), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n800), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n796), .B(new_n611), .C1(new_n807), .C2(KEYINPUT55), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n802), .A2(new_n801), .A3(new_n628), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT114), .B1(new_n804), .B2(new_n805), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT55), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n629), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n676), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n815));
  INV_X1    g614(.A(new_n793), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n789), .A2(new_n792), .B1(new_n533), .B2(new_n534), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n541), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n536), .B2(new_n675), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n815), .A2(new_n813), .B1(new_n632), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n814), .B1(new_n820), .B2(new_n612), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n786), .B1(new_n821), .B2(new_n673), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n694), .A2(new_n459), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n456), .A2(new_n447), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n304), .A3(new_n543), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n630), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n828), .A2(new_n611), .A3(new_n831), .A4(new_n796), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n632), .A2(new_n819), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n543), .B1(new_n829), .B2(new_n830), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n828), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n835), .B2(new_n611), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n785), .B1(new_n836), .B2(new_n674), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n456), .A3(new_n495), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n457), .A3(new_n676), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n827), .B1(new_n839), .B2(new_n304), .ZN(G1340gat));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n823), .A3(new_n633), .A4(new_n825), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n841), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT116), .B1(new_n841), .B2(G120gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n838), .A2(new_n457), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n633), .A2(new_n286), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT117), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n842), .A2(new_n843), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT118), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n826), .B2(new_n674), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n575), .A2(new_n291), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT119), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n612), .A2(new_n447), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n293), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n826), .B2(new_n612), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n837), .B2(new_n281), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n786), .B1(new_n821), .B2(new_n575), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n459), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT120), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT57), .A4(new_n459), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n493), .A2(new_n825), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n676), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n493), .A2(new_n459), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n822), .A2(new_n545), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n457), .ZN(new_n871));
  INV_X1    g670(.A(G141gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n676), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(G148gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT59), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n632), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n633), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n837), .A2(new_n859), .A3(new_n281), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n861), .B2(new_n459), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G148gat), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT121), .B1(new_n888), .B2(KEYINPUT59), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n785), .B1(new_n836), .B2(new_n574), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n859), .B1(new_n890), .B2(new_n281), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n459), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n883), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n893), .C2(new_n879), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n882), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n879), .A3(new_n633), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1345gat));
  OAI21_X1  g697(.A(G155gat), .B1(new_n881), .B2(new_n674), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n871), .A2(new_n246), .A3(new_n575), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1346gat));
  NAND4_X1  g700(.A1(new_n863), .A2(new_n611), .A3(new_n865), .A4(new_n866), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G162gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n870), .A2(new_n247), .A3(new_n853), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(KEYINPUT122), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n495), .A2(new_n457), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT124), .Z(new_n911));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n837), .B2(new_n545), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n822), .A2(KEYINPUT123), .A3(new_n456), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n676), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n545), .A2(new_n457), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n824), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(G169gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(new_n543), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n916), .A2(new_n920), .ZN(G1348gat));
  INV_X1    g720(.A(G176gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n915), .A2(new_n922), .A3(new_n633), .ZN(new_n923));
  OAI21_X1  g722(.A(G176gat), .B1(new_n918), .B2(new_n632), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1349gat));
  OAI21_X1  g724(.A(G183gat), .B1(new_n918), .B2(new_n674), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n575), .A2(new_n380), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n915), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n915), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n915), .A2(new_n356), .A3(new_n611), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n824), .A2(new_n611), .A3(new_n917), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(G190gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n937), .B2(G190gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n913), .A2(new_n914), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n869), .A2(new_n447), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT126), .B(G197gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n676), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n891), .A2(new_n892), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n493), .A3(new_n917), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n543), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n950), .B2(new_n946), .ZN(G1352gat));
  NOR2_X1   g750(.A1(new_n632), .A2(G204gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n945), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT127), .B1(new_n949), .B2(new_n632), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n949), .A2(KEYINPUT127), .A3(new_n632), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n954), .B(new_n956), .C1(new_n958), .C2(new_n959), .ZN(G1353gat));
  NAND4_X1  g759(.A1(new_n945), .A2(new_n212), .A3(new_n213), .A4(new_n575), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n948), .A2(new_n493), .A3(new_n575), .A4(new_n917), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n949), .B2(new_n612), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n611), .A2(new_n211), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n944), .B2(new_n967), .ZN(G1355gat));
endmodule


