

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802;

  NOR2_X1 U383 ( .A1(n634), .A2(n633), .ZN(n644) );
  OR2_X1 U384 ( .A1(n445), .A2(n443), .ZN(n612) );
  NAND2_X2 U385 ( .A1(n406), .A2(n391), .ZN(n656) );
  AND2_X2 U386 ( .A1(n390), .A2(n405), .ZN(n406) );
  XNOR2_X2 U387 ( .A(n452), .B(KEYINPUT104), .ZN(n674) );
  XNOR2_X2 U388 ( .A(n511), .B(n510), .ZN(n530) );
  XNOR2_X2 U389 ( .A(n468), .B(G128), .ZN(n511) );
  XNOR2_X2 U390 ( .A(n620), .B(KEYINPUT40), .ZN(n800) );
  AND2_X2 U391 ( .A1(n648), .A2(n764), .ZN(n620) );
  NOR2_X1 U392 ( .A1(n378), .A2(n675), .ZN(n679) );
  AND2_X1 U393 ( .A1(n424), .A2(n420), .ZN(n419) );
  NAND2_X1 U394 ( .A1(n383), .A2(n379), .ZN(n797) );
  NOR2_X1 U395 ( .A1(n628), .A2(n409), .ZN(n408) );
  AND2_X1 U396 ( .A1(n459), .A2(n373), .ZN(n457) );
  AND2_X1 U397 ( .A1(n441), .A2(n440), .ZN(n439) );
  AND2_X1 U398 ( .A1(n651), .A2(KEYINPUT82), .ZN(n404) );
  XNOR2_X1 U399 ( .A(n787), .B(n531), .ZN(n543) );
  XNOR2_X1 U400 ( .A(n465), .B(KEYINPUT3), .ZN(n427) );
  BUF_X2 U401 ( .A(n701), .Z(n791) );
  XNOR2_X2 U402 ( .A(n393), .B(n365), .ZN(n614) );
  NAND2_X2 U403 ( .A1(n389), .A2(n399), .ZN(n393) );
  XNOR2_X2 U404 ( .A(n534), .B(n464), .ZN(n428) );
  XNOR2_X2 U405 ( .A(n775), .B(n473), .ZN(n665) );
  XNOR2_X2 U406 ( .A(n428), .B(n541), .ZN(n775) );
  NAND2_X1 U407 ( .A1(n695), .A2(n693), .ZN(n447) );
  XNOR2_X1 U408 ( .A(n530), .B(n529), .ZN(n787) );
  XNOR2_X1 U409 ( .A(G137), .B(KEYINPUT4), .ZN(n528) );
  XNOR2_X1 U410 ( .A(G146), .B(G125), .ZN(n494) );
  NAND2_X1 U411 ( .A1(n401), .A2(n652), .ZN(n400) );
  INV_X1 U412 ( .A(n478), .ZN(n401) );
  NAND2_X1 U413 ( .A1(n447), .A2(n446), .ZN(n445) );
  NAND2_X1 U414 ( .A1(G469), .A2(n556), .ZN(n444) );
  XNOR2_X1 U415 ( .A(G119), .B(G116), .ZN(n431) );
  AND2_X1 U416 ( .A1(n388), .A2(n387), .ZN(n398) );
  XNOR2_X1 U417 ( .A(n583), .B(KEYINPUT107), .ZN(n388) );
  INV_X1 U418 ( .A(KEYINPUT86), .ZN(n450) );
  INV_X1 U419 ( .A(KEYINPUT85), .ZN(n415) );
  INV_X1 U420 ( .A(KEYINPUT101), .ZN(n497) );
  XNOR2_X1 U421 ( .A(G113), .B(G122), .ZN(n502) );
  XOR2_X1 U422 ( .A(KEYINPUT11), .B(G104), .Z(n503) );
  INV_X1 U423 ( .A(KEYINPUT109), .ZN(n411) );
  NAND2_X1 U424 ( .A1(n650), .A2(n478), .ZN(n402) );
  XNOR2_X1 U425 ( .A(n509), .B(n508), .ZN(n588) );
  NOR2_X1 U426 ( .A1(G902), .A2(n657), .ZN(n509) );
  NOR2_X1 U427 ( .A1(G953), .A2(G237), .ZN(n537) );
  INV_X1 U428 ( .A(KEYINPUT10), .ZN(n492) );
  INV_X1 U429 ( .A(G146), .ZN(n531) );
  INV_X1 U430 ( .A(KEYINPUT79), .ZN(n433) );
  NOR2_X1 U431 ( .A1(n363), .A2(n386), .ZN(n385) );
  NAND2_X1 U432 ( .A1(n439), .A2(n438), .ZN(n386) );
  NAND2_X1 U433 ( .A1(n435), .A2(n434), .ZN(n384) );
  INV_X1 U434 ( .A(n442), .ZN(n434) );
  NAND2_X1 U435 ( .A1(n364), .A2(n382), .ZN(n381) );
  NAND2_X1 U436 ( .A1(n743), .A2(n439), .ZN(n382) );
  NAND2_X1 U437 ( .A1(n439), .A2(n442), .ZN(n437) );
  XNOR2_X1 U438 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n526) );
  INV_X1 U439 ( .A(KEYINPUT77), .ZN(n397) );
  INV_X2 U440 ( .A(G953), .ZN(n793) );
  NOR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n476) );
  XOR2_X1 U442 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n496) );
  XNOR2_X1 U443 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n495) );
  XNOR2_X1 U444 ( .A(G143), .B(G131), .ZN(n498) );
  XNOR2_X1 U445 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n474) );
  NOR2_X1 U446 ( .A1(n423), .A2(n422), .ZN(n421) );
  NAND2_X1 U447 ( .A1(n693), .A2(G902), .ZN(n446) );
  XNOR2_X1 U448 ( .A(n516), .B(n515), .ZN(n547) );
  XNOR2_X1 U449 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n515) );
  NAND2_X1 U450 ( .A1(n392), .A2(n651), .ZN(n405) );
  NAND2_X1 U451 ( .A1(n652), .A2(KEYINPUT82), .ZN(n454) );
  INV_X1 U452 ( .A(G143), .ZN(n468) );
  XNOR2_X1 U453 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n470) );
  NOR2_X1 U454 ( .A1(n706), .A2(KEYINPUT2), .ZN(n700) );
  INV_X1 U455 ( .A(n630), .ZN(n387) );
  NAND2_X1 U456 ( .A1(n573), .A2(n436), .ZN(n442) );
  INV_X1 U457 ( .A(n604), .ZN(n440) );
  XOR2_X1 U458 ( .A(G101), .B(KEYINPUT5), .Z(n539) );
  XNOR2_X1 U459 ( .A(G128), .B(G137), .ZN(n549) );
  INV_X1 U460 ( .A(G134), .ZN(n510) );
  XNOR2_X1 U461 ( .A(G116), .B(G122), .ZN(n512) );
  XOR2_X1 U462 ( .A(KEYINPUT102), .B(G107), .Z(n513) );
  XNOR2_X1 U463 ( .A(n507), .B(n506), .ZN(n657) );
  XNOR2_X1 U464 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U465 ( .A(n412), .B(n410), .ZN(n613) );
  XNOR2_X1 U466 ( .A(n611), .B(n411), .ZN(n410) );
  NOR2_X1 U467 ( .A1(n714), .A2(n713), .ZN(n623) );
  AND2_X1 U468 ( .A1(n602), .A2(n395), .ZN(n394) );
  INV_X1 U469 ( .A(n634), .ZN(n395) );
  AND2_X1 U470 ( .A1(n545), .A2(n546), .ZN(n460) );
  OR2_X1 U471 ( .A1(n545), .A2(n546), .ZN(n458) );
  XOR2_X1 U472 ( .A(n521), .B(G478), .Z(n589) );
  INV_X1 U473 ( .A(n588), .ZN(n590) );
  XNOR2_X1 U474 ( .A(KEYINPUT16), .B(G122), .ZN(n464) );
  XNOR2_X1 U475 ( .A(n543), .B(n535), .ZN(n695) );
  XNOR2_X1 U476 ( .A(n705), .B(n433), .ZN(n432) );
  AND2_X1 U477 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U478 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X1 U479 ( .A(n568), .B(n567), .ZN(n672) );
  NOR2_X1 U480 ( .A1(n590), .A2(n589), .ZN(n764) );
  AND2_X1 U481 ( .A1(n743), .A2(KEYINPUT34), .ZN(n363) );
  AND2_X1 U482 ( .A1(n437), .A2(n376), .ZN(n364) );
  XNOR2_X1 U483 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n365) );
  NAND2_X1 U484 ( .A1(n416), .A2(n419), .ZN(n706) );
  INV_X1 U485 ( .A(n570), .ZN(n727) );
  XOR2_X1 U486 ( .A(n536), .B(KEYINPUT1), .Z(n367) );
  AND2_X1 U487 ( .A1(n618), .A2(n617), .ZN(n368) );
  XOR2_X1 U488 ( .A(KEYINPUT30), .B(n601), .Z(n369) );
  AND2_X1 U489 ( .A1(n416), .A2(n404), .ZN(n370) );
  AND2_X1 U490 ( .A1(n369), .A2(n394), .ZN(n371) );
  AND2_X1 U491 ( .A1(n399), .A2(n402), .ZN(n372) );
  AND2_X1 U492 ( .A1(n458), .A2(n562), .ZN(n373) );
  AND2_X1 U493 ( .A1(n402), .A2(n710), .ZN(n374) );
  XOR2_X1 U494 ( .A(n490), .B(KEYINPUT0), .Z(n375) );
  XOR2_X1 U495 ( .A(KEYINPUT83), .B(KEYINPUT35), .Z(n376) );
  NOR2_X1 U496 ( .A1(n438), .A2(n436), .ZN(n377) );
  INV_X1 U497 ( .A(KEYINPUT45), .ZN(n422) );
  XNOR2_X1 U498 ( .A(n656), .B(KEYINPUT64), .ZN(n378) );
  XNOR2_X1 U499 ( .A(n656), .B(KEYINPUT64), .ZN(n692) );
  NAND2_X1 U500 ( .A1(n614), .A2(n489), .ZN(n491) );
  NAND2_X1 U501 ( .A1(n743), .A2(n377), .ZN(n380) );
  NAND2_X1 U502 ( .A1(n570), .A2(n569), .ZN(n583) );
  XNOR2_X2 U503 ( .A(n612), .B(n367), .ZN(n570) );
  OR2_X1 U504 ( .A1(n665), .A2(n400), .ZN(n399) );
  AND2_X2 U505 ( .A1(n403), .A2(n374), .ZN(n389) );
  XNOR2_X1 U506 ( .A(n581), .B(n582), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n453), .A2(n722), .ZN(n452) );
  XOR2_X2 U508 ( .A(KEYINPUT6), .B(n725), .Z(n630) );
  NAND2_X1 U509 ( .A1(n370), .A2(n419), .ZN(n390) );
  NAND2_X1 U510 ( .A1(n655), .A2(n706), .ZN(n391) );
  NAND2_X1 U511 ( .A1(n707), .A2(n454), .ZN(n392) );
  NAND2_X1 U512 ( .A1(n564), .A2(n396), .ZN(n565) );
  XNOR2_X1 U513 ( .A(n630), .B(n397), .ZN(n396) );
  XNOR2_X1 U514 ( .A(n426), .B(n415), .ZN(n425) );
  XNOR2_X2 U515 ( .A(n398), .B(n571), .ZN(n743) );
  XNOR2_X1 U516 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U517 ( .A1(n403), .A2(n372), .ZN(n603) );
  NAND2_X1 U518 ( .A1(n665), .A2(n478), .ZN(n403) );
  NAND2_X1 U519 ( .A1(n407), .A2(n649), .ZN(n701) );
  XNOR2_X1 U520 ( .A(n408), .B(KEYINPUT48), .ZN(n407) );
  NAND2_X1 U521 ( .A1(n643), .A2(n368), .ZN(n409) );
  NAND2_X1 U522 ( .A1(n610), .A2(n413), .ZN(n412) );
  NOR2_X1 U523 ( .A1(n725), .A2(n634), .ZN(n413) );
  NAND2_X1 U524 ( .A1(n414), .A2(n421), .ZN(n420) );
  NAND2_X1 U525 ( .A1(n414), .A2(n579), .ZN(n417) );
  NAND2_X1 U526 ( .A1(n575), .A2(n574), .ZN(n414) );
  NOR2_X1 U527 ( .A1(n425), .A2(KEYINPUT45), .ZN(n418) );
  NAND2_X1 U528 ( .A1(n418), .A2(n417), .ZN(n416) );
  INV_X1 U529 ( .A(n579), .ZN(n423) );
  NAND2_X1 U530 ( .A1(n425), .A2(KEYINPUT45), .ZN(n424) );
  NAND2_X1 U531 ( .A1(n594), .A2(n595), .ZN(n426) );
  XNOR2_X2 U532 ( .A(n427), .B(n431), .ZN(n541) );
  XNOR2_X2 U533 ( .A(n430), .B(n429), .ZN(n534) );
  XNOR2_X2 U534 ( .A(G110), .B(G107), .ZN(n429) );
  XNOR2_X2 U535 ( .A(G104), .B(G101), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n578), .B(n450), .ZN(n449) );
  NOR2_X1 U537 ( .A1(n432), .A2(n709), .ZN(n748) );
  NAND2_X2 U538 ( .A1(n457), .A2(n455), .ZN(n673) );
  NAND2_X1 U539 ( .A1(n449), .A2(n451), .ZN(n448) );
  INV_X1 U540 ( .A(n743), .ZN(n435) );
  NAND2_X1 U541 ( .A1(n586), .A2(KEYINPUT34), .ZN(n441) );
  INV_X1 U542 ( .A(KEYINPUT34), .ZN(n436) );
  INV_X1 U543 ( .A(n376), .ZN(n438) );
  NOR2_X1 U544 ( .A1(n695), .A2(n444), .ZN(n443) );
  OR2_X2 U545 ( .A1(n677), .A2(G902), .ZN(n544) );
  XNOR2_X1 U546 ( .A(n448), .B(n576), .ZN(n575) );
  INV_X1 U547 ( .A(n797), .ZN(n451) );
  NAND2_X1 U548 ( .A1(n673), .A2(n672), .ZN(n578) );
  XNOR2_X1 U549 ( .A(n580), .B(KEYINPUT106), .ZN(n461) );
  NOR2_X2 U550 ( .A1(n563), .A2(n570), .ZN(n580) );
  NAND2_X1 U551 ( .A1(n674), .A2(n592), .ZN(n593) );
  INV_X1 U552 ( .A(n706), .ZN(n366) );
  NAND2_X1 U553 ( .A1(n456), .A2(KEYINPUT66), .ZN(n455) );
  INV_X1 U554 ( .A(n461), .ZN(n456) );
  NAND2_X1 U555 ( .A1(n461), .A2(n460), .ZN(n459) );
  BUF_X1 U556 ( .A(n682), .Z(n688) );
  XOR2_X1 U557 ( .A(n548), .B(n785), .Z(n462) );
  AND2_X1 U558 ( .A1(n642), .A2(KEYINPUT47), .ZN(n463) );
  INV_X1 U559 ( .A(KEYINPUT46), .ZN(n626) );
  NOR2_X1 U560 ( .A1(n801), .A2(n463), .ZN(n643) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U563 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n571) );
  INV_X1 U564 ( .A(n726), .ZN(n569) );
  INV_X1 U565 ( .A(KEYINPUT66), .ZN(n546) );
  NAND2_X1 U566 ( .A1(n688), .A2(G217), .ZN(n685) );
  XNOR2_X1 U567 ( .A(n685), .B(n684), .ZN(n687) );
  XNOR2_X2 U568 ( .A(G113), .B(KEYINPUT70), .ZN(n465) );
  XNOR2_X1 U569 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n467) );
  NAND2_X1 U570 ( .A1(n793), .A2(G224), .ZN(n466) );
  XNOR2_X1 U571 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U572 ( .A(n511), .B(n469), .ZN(n472) );
  XNOR2_X1 U573 ( .A(n494), .B(n470), .ZN(n471) );
  XNOR2_X1 U574 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U575 ( .A(n474), .B(G902), .ZN(n652) );
  INV_X1 U576 ( .A(n652), .ZN(n650) );
  INV_X1 U577 ( .A(KEYINPUT75), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n480) );
  INV_X1 U579 ( .A(n480), .ZN(n477) );
  NAND2_X1 U580 ( .A1(n477), .A2(G210), .ZN(n478) );
  INV_X1 U581 ( .A(G214), .ZN(n479) );
  OR2_X1 U582 ( .A1(n480), .A2(n479), .ZN(n710) );
  NAND2_X1 U583 ( .A1(G234), .A2(G237), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n481), .B(KEYINPUT14), .ZN(n482) );
  XNOR2_X1 U585 ( .A(KEYINPUT74), .B(n482), .ZN(n486) );
  NAND2_X1 U586 ( .A1(n486), .A2(G902), .ZN(n483) );
  XNOR2_X1 U587 ( .A(KEYINPUT94), .B(n483), .ZN(n596) );
  XOR2_X1 U588 ( .A(G898), .B(KEYINPUT92), .Z(n780) );
  NAND2_X1 U589 ( .A1(n780), .A2(G953), .ZN(n484) );
  XOR2_X1 U590 ( .A(KEYINPUT93), .B(n484), .Z(n776) );
  NOR2_X1 U591 ( .A1(n596), .A2(n776), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n485), .B(KEYINPUT95), .ZN(n488) );
  NAND2_X1 U593 ( .A1(G952), .A2(n486), .ZN(n738) );
  NOR2_X1 U594 ( .A1(n738), .A2(G953), .ZN(n599) );
  INV_X1 U595 ( .A(n599), .ZN(n487) );
  NAND2_X1 U596 ( .A1(n488), .A2(n487), .ZN(n489) );
  INV_X1 U597 ( .A(KEYINPUT87), .ZN(n490) );
  XNOR2_X2 U598 ( .A(n491), .B(n375), .ZN(n572) );
  XNOR2_X1 U599 ( .A(n492), .B(G140), .ZN(n493) );
  XNOR2_X1 U600 ( .A(n494), .B(n493), .ZN(n785) );
  XNOR2_X1 U601 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n501), .B(n785), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n505) );
  AND2_X1 U604 ( .A1(G214), .A2(n537), .ZN(n504) );
  XNOR2_X1 U605 ( .A(KEYINPUT13), .B(G475), .ZN(n508) );
  XNOR2_X1 U606 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U607 ( .A(n530), .B(n514), .ZN(n520) );
  NAND2_X1 U608 ( .A1(n793), .A2(G234), .ZN(n516) );
  NAND2_X1 U609 ( .A1(G217), .A2(n547), .ZN(n518) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n517) );
  XNOR2_X1 U611 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n519), .B(n520), .ZN(n689) );
  NOR2_X1 U613 ( .A1(n689), .A2(G902), .ZN(n521) );
  NOR2_X1 U614 ( .A1(n588), .A2(n589), .ZN(n621) );
  NAND2_X1 U615 ( .A1(n652), .A2(G234), .ZN(n522) );
  XNOR2_X1 U616 ( .A(KEYINPUT20), .B(n522), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n557), .A2(G221), .ZN(n523) );
  XNOR2_X1 U618 ( .A(KEYINPUT21), .B(n523), .ZN(n609) );
  INV_X1 U619 ( .A(n609), .ZN(n721) );
  NAND2_X1 U620 ( .A1(n621), .A2(n721), .ZN(n524) );
  XNOR2_X1 U621 ( .A(n524), .B(KEYINPUT103), .ZN(n525) );
  NAND2_X1 U622 ( .A1(n572), .A2(n525), .ZN(n527) );
  XNOR2_X1 U623 ( .A(n527), .B(n526), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n528), .B(G131), .ZN(n529) );
  NAND2_X1 U625 ( .A1(G227), .A2(n793), .ZN(n532) );
  XNOR2_X1 U626 ( .A(n532), .B(G140), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n534), .B(n533), .ZN(n535) );
  INV_X1 U628 ( .A(G469), .ZN(n693) );
  INV_X1 U629 ( .A(KEYINPUT67), .ZN(n536) );
  NAND2_X1 U630 ( .A1(n537), .A2(G210), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U633 ( .A(n543), .B(n542), .ZN(n677) );
  INV_X1 U634 ( .A(G472), .ZN(n675) );
  XNOR2_X2 U635 ( .A(n544), .B(n675), .ZN(n725) );
  INV_X1 U636 ( .A(n725), .ZN(n600) );
  INV_X1 U637 ( .A(n600), .ZN(n545) );
  NAND2_X1 U638 ( .A1(G221), .A2(n547), .ZN(n548) );
  XOR2_X1 U639 ( .A(G110), .B(G119), .Z(n550) );
  XNOR2_X1 U640 ( .A(n550), .B(n549), .ZN(n554) );
  XOR2_X1 U641 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n552) );
  XNOR2_X1 U642 ( .A(KEYINPUT24), .B(KEYINPUT76), .ZN(n551) );
  XNOR2_X1 U643 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U644 ( .A(n554), .B(n553), .Z(n555) );
  XNOR2_X1 U645 ( .A(n462), .B(n555), .ZN(n683) );
  INV_X1 U646 ( .A(G902), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n683), .A2(n556), .ZN(n561) );
  NAND2_X1 U648 ( .A1(G217), .A2(n557), .ZN(n559) );
  INV_X1 U649 ( .A(KEYINPUT25), .ZN(n558) );
  XNOR2_X1 U650 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X2 U651 ( .A(n561), .B(n560), .ZN(n722) );
  INV_X1 U652 ( .A(n722), .ZN(n562) );
  BUF_X1 U653 ( .A(n563), .Z(n566) );
  NOR2_X1 U654 ( .A1(n727), .A2(n722), .ZN(n564) );
  NOR2_X1 U655 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U656 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n567) );
  NAND2_X1 U657 ( .A1(n721), .A2(n722), .ZN(n726) );
  BUF_X1 U658 ( .A(n572), .Z(n573) );
  INV_X1 U659 ( .A(n573), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n588), .A2(n589), .ZN(n604) );
  INV_X1 U661 ( .A(KEYINPUT44), .ZN(n574) );
  INV_X1 U662 ( .A(KEYINPUT71), .ZN(n576) );
  NAND2_X1 U663 ( .A1(n576), .A2(KEYINPUT44), .ZN(n577) );
  OR2_X1 U664 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U665 ( .A1(n797), .A2(KEYINPUT44), .ZN(n595) );
  INV_X1 U666 ( .A(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U667 ( .A1(n580), .A2(n630), .ZN(n581) );
  NOR2_X1 U668 ( .A1(n583), .A2(n725), .ZN(n732) );
  NAND2_X1 U669 ( .A1(n732), .A2(n573), .ZN(n585) );
  XNOR2_X1 U670 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n584) );
  XNOR2_X1 U671 ( .A(n585), .B(n584), .ZN(n770) );
  NOR2_X1 U672 ( .A1(n612), .A2(n726), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n602), .A2(n545), .ZN(n587) );
  OR2_X1 U674 ( .A1(n587), .A2(n586), .ZN(n753) );
  NAND2_X1 U675 ( .A1(n770), .A2(n753), .ZN(n591) );
  INV_X1 U676 ( .A(n764), .ZN(n767) );
  NAND2_X1 U677 ( .A1(n590), .A2(n589), .ZN(n771) );
  NAND2_X1 U678 ( .A1(n767), .A2(n771), .ZN(n640) );
  NAND2_X1 U679 ( .A1(n591), .A2(n640), .ZN(n592) );
  XNOR2_X1 U680 ( .A(n593), .B(KEYINPUT105), .ZN(n594) );
  OR2_X1 U681 ( .A1(n793), .A2(n596), .ZN(n597) );
  NOR2_X1 U682 ( .A1(G900), .A2(n597), .ZN(n598) );
  NOR2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n634) );
  NAND2_X1 U684 ( .A1(n600), .A2(n710), .ZN(n601) );
  NOR2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n605) );
  AND2_X1 U686 ( .A1(n371), .A2(n605), .ZN(n762) );
  NOR2_X1 U687 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n606) );
  NOR2_X1 U688 ( .A1(n762), .A2(n606), .ZN(n618) );
  INV_X1 U689 ( .A(n640), .ZN(n715) );
  NOR2_X1 U690 ( .A1(n715), .A2(KEYINPUT47), .ZN(n607) );
  XNOR2_X1 U691 ( .A(n607), .B(KEYINPUT73), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n608), .A2(KEYINPUT80), .ZN(n616) );
  XNOR2_X1 U693 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n611) );
  NOR2_X1 U694 ( .A1(n722), .A2(n609), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n624), .A2(n614), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(KEYINPUT78), .ZN(n639) );
  INV_X1 U698 ( .A(n639), .ZN(n765) );
  NAND2_X1 U699 ( .A1(n616), .A2(n765), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n603), .B(KEYINPUT38), .ZN(n711) );
  NAND2_X1 U701 ( .A1(n371), .A2(n711), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT39), .ZN(n648) );
  NAND2_X1 U703 ( .A1(n711), .A2(n710), .ZN(n714) );
  INV_X1 U704 ( .A(n621), .ZN(n713) );
  XNOR2_X1 U705 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n622) );
  XNOR2_X1 U706 ( .A(n623), .B(n622), .ZN(n741) );
  NAND2_X1 U707 ( .A1(n741), .A2(n624), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT42), .B(n625), .Z(n798) );
  NOR2_X1 U709 ( .A1(n800), .A2(n798), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n710), .A2(n721), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n767), .A2(n629), .ZN(n632) );
  NOR2_X1 U712 ( .A1(n722), .A2(n630), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  INV_X1 U714 ( .A(n603), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n644), .A2(n635), .ZN(n636) );
  XNOR2_X1 U716 ( .A(n636), .B(KEYINPUT36), .ZN(n637) );
  NOR2_X1 U717 ( .A1(n637), .A2(n727), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n638), .B(KEYINPUT112), .ZN(n801) );
  NAND2_X1 U719 ( .A1(n639), .A2(KEYINPUT80), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U721 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n646) );
  NAND2_X1 U722 ( .A1(n644), .A2(n727), .ZN(n645) );
  XOR2_X1 U723 ( .A(n646), .B(n645), .Z(n647) );
  NAND2_X1 U724 ( .A1(n647), .A2(n603), .ZN(n671) );
  INV_X1 U725 ( .A(n771), .ZN(n759) );
  NAND2_X1 U726 ( .A1(n648), .A2(n759), .ZN(n774) );
  AND2_X1 U727 ( .A1(n671), .A2(n774), .ZN(n649) );
  INV_X1 U728 ( .A(n701), .ZN(n707) );
  NAND2_X1 U729 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  NOR2_X1 U730 ( .A1(n652), .A2(KEYINPUT82), .ZN(n653) );
  NOR2_X1 U731 ( .A1(n653), .A2(KEYINPUT2), .ZN(n654) );
  NOR2_X1 U732 ( .A1(n791), .A2(n654), .ZN(n655) );
  INV_X1 U733 ( .A(n692), .ZN(n682) );
  NAND2_X1 U734 ( .A1(n682), .A2(G475), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n657), .B(KEYINPUT59), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n661) );
  NOR2_X1 U737 ( .A1(n793), .A2(G952), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(KEYINPUT89), .ZN(n686) );
  NAND2_X1 U739 ( .A1(n661), .A2(n686), .ZN(n663) );
  INV_X1 U740 ( .A(KEYINPUT60), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(G60) );
  NAND2_X1 U742 ( .A1(n682), .A2(G210), .ZN(n667) );
  XNOR2_X1 U743 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n668), .A2(n686), .ZN(n670) );
  INV_X1 U747 ( .A(KEYINPUT56), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(G51) );
  XNOR2_X1 U749 ( .A(n671), .B(G140), .ZN(G42) );
  XNOR2_X1 U750 ( .A(n672), .B(G119), .ZN(G21) );
  XNOR2_X1 U751 ( .A(n673), .B(G110), .ZN(G12) );
  XNOR2_X1 U752 ( .A(n674), .B(G101), .ZN(G3) );
  XOR2_X1 U753 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n676) );
  XNOR2_X1 U754 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U755 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U756 ( .A1(n680), .A2(n686), .ZN(n681) );
  XNOR2_X1 U757 ( .A(n681), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U758 ( .A(n683), .ZN(n684) );
  INV_X1 U759 ( .A(n686), .ZN(n698) );
  NOR2_X1 U760 ( .A1(n687), .A2(n698), .ZN(G66) );
  NAND2_X1 U761 ( .A1(n688), .A2(G478), .ZN(n690) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n691), .A2(n698), .ZN(G63) );
  NOR2_X1 U764 ( .A1(n378), .A2(n693), .ZN(n697) );
  XNOR2_X1 U765 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(G54) );
  XNOR2_X1 U769 ( .A(n700), .B(KEYINPUT81), .ZN(n704) );
  INV_X1 U770 ( .A(KEYINPUT2), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n791), .A2(n702), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n707), .A2(KEYINPUT2), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n366), .A2(n708), .ZN(n709) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U779 ( .A(n718), .B(KEYINPUT120), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n743), .A2(n719), .ZN(n720) );
  XNOR2_X1 U781 ( .A(n720), .B(KEYINPUT121), .ZN(n736) );
  NOR2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U783 ( .A(n723), .B(KEYINPUT49), .ZN(n724) );
  NAND2_X1 U784 ( .A1(n725), .A2(n724), .ZN(n730) );
  NAND2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U786 ( .A(KEYINPUT50), .B(n728), .Z(n729) );
  NOR2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U788 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U789 ( .A(KEYINPUT51), .B(n733), .ZN(n734) );
  NAND2_X1 U790 ( .A1(n734), .A2(n741), .ZN(n735) );
  NAND2_X1 U791 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U792 ( .A(KEYINPUT52), .B(n737), .Z(n739) );
  NOR2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U794 ( .A(KEYINPUT122), .B(n740), .Z(n746) );
  INV_X1 U795 ( .A(n741), .ZN(n742) );
  NOR2_X1 U796 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U797 ( .A1(n744), .A2(G953), .ZN(n745) );
  NAND2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U799 ( .A1(n748), .A2(n747), .ZN(n750) );
  XOR2_X1 U800 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(G75) );
  NOR2_X1 U802 ( .A1(n753), .A2(n767), .ZN(n751) );
  XOR2_X1 U803 ( .A(KEYINPUT114), .B(n751), .Z(n752) );
  XNOR2_X1 U804 ( .A(G104), .B(n752), .ZN(G6) );
  NOR2_X1 U805 ( .A1(n753), .A2(n771), .ZN(n758) );
  XOR2_X1 U806 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n755) );
  XNOR2_X1 U807 ( .A(G107), .B(KEYINPUT115), .ZN(n754) );
  XNOR2_X1 U808 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U809 ( .A(KEYINPUT26), .B(n756), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n758), .B(n757), .ZN(G9) );
  XOR2_X1 U811 ( .A(G128), .B(KEYINPUT29), .Z(n761) );
  NAND2_X1 U812 ( .A1(n759), .A2(n765), .ZN(n760) );
  XNOR2_X1 U813 ( .A(n761), .B(n760), .ZN(G30) );
  XNOR2_X1 U814 ( .A(G143), .B(n762), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n763), .B(KEYINPUT117), .ZN(G45) );
  NAND2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n766), .B(G146), .ZN(G48) );
  NOR2_X1 U818 ( .A1(n767), .A2(n770), .ZN(n768) );
  XOR2_X1 U819 ( .A(KEYINPUT118), .B(n768), .Z(n769) );
  XNOR2_X1 U820 ( .A(G113), .B(n769), .ZN(G15) );
  NOR2_X1 U821 ( .A1(n771), .A2(n770), .ZN(n773) );
  XNOR2_X1 U822 ( .A(G116), .B(KEYINPUT119), .ZN(n772) );
  XNOR2_X1 U823 ( .A(n773), .B(n772), .ZN(G18) );
  XNOR2_X1 U824 ( .A(G134), .B(n774), .ZN(G36) );
  XOR2_X1 U825 ( .A(KEYINPUT124), .B(n775), .Z(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n784) );
  NOR2_X1 U827 ( .A1(n366), .A2(G953), .ZN(n782) );
  NAND2_X1 U828 ( .A1(G953), .A2(G224), .ZN(n778) );
  XOR2_X1 U829 ( .A(KEYINPUT61), .B(n778), .Z(n779) );
  NOR2_X1 U830 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U832 ( .A(n784), .B(n783), .ZN(G69) );
  XOR2_X1 U833 ( .A(n785), .B(KEYINPUT125), .Z(n786) );
  XOR2_X1 U834 ( .A(n787), .B(n786), .Z(n792) );
  XOR2_X1 U835 ( .A(n792), .B(KEYINPUT126), .Z(n788) );
  XNOR2_X1 U836 ( .A(G227), .B(n788), .ZN(n789) );
  NAND2_X1 U837 ( .A1(G900), .A2(n789), .ZN(n790) );
  NAND2_X1 U838 ( .A1(n790), .A2(G953), .ZN(n796) );
  XOR2_X1 U839 ( .A(n792), .B(n791), .Z(n794) );
  NAND2_X1 U840 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U841 ( .A1(n796), .A2(n795), .ZN(G72) );
  XOR2_X1 U842 ( .A(n797), .B(G122), .Z(G24) );
  XNOR2_X1 U843 ( .A(G137), .B(KEYINPUT127), .ZN(n799) );
  XNOR2_X1 U844 ( .A(n799), .B(n798), .ZN(G39) );
  XOR2_X1 U845 ( .A(n800), .B(G131), .Z(G33) );
  XNOR2_X1 U846 ( .A(G125), .B(KEYINPUT37), .ZN(n802) );
  XNOR2_X1 U847 ( .A(n802), .B(n801), .ZN(G27) );
endmodule

