//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(G113), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(KEYINPUT69), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n464), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(new_n470), .A3(KEYINPUT3), .A4(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n463), .B2(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  AND2_X1   g053(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n474), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n475), .A3(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n460), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n475), .A2(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n474), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n474), .A2(G126), .A3(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n494), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n506), .B1(new_n502), .B2(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  XOR2_X1   g089(.A(KEYINPUT73), .B(G88), .Z(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G50), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n503), .A2(new_n506), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n502), .A2(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(new_n513), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n511), .A2(KEYINPUT75), .A3(new_n512), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(G543), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n523), .B1(new_n526), .B2(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n521), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n509), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n531), .A2(new_n537), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n507), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n509), .B1(new_n544), .B2(KEYINPUT76), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(KEYINPUT76), .B2(new_n544), .ZN(new_n546));
  INV_X1    g121(.A(new_n531), .ZN(new_n547));
  INV_X1    g122(.A(new_n526), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n547), .A2(G43), .B1(new_n548), .B2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G860), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  AOI21_X1  g132(.A(new_n505), .B1(new_n513), .B2(new_n528), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n558), .A2(G53), .A3(new_n530), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n526), .A2(KEYINPUT78), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n507), .A2(new_n562), .A3(new_n513), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(KEYINPUT79), .B(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n542), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n560), .A2(new_n565), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n574));
  INV_X1    g149(.A(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n531), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n558), .A2(KEYINPUT80), .A3(G49), .A4(new_n530), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n561), .A2(G87), .A3(new_n563), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n583), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n561), .A2(G86), .A3(new_n563), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n547), .A2(G47), .B1(new_n548), .B2(G85), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n509), .B2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n564), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n507), .A2(G66), .ZN(new_n596));
  INV_X1    g171(.A(G79), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT81), .B1(new_n597), .B2(new_n505), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n597), .A2(new_n505), .A3(KEYINPUT81), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(new_n547), .B2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n592), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n592), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  OR3_X1    g181(.A1(G168), .A2(KEYINPUT82), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT82), .B1(G168), .B2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n606), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(G297));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(G280));
  AOI21_X1  g186(.A(new_n602), .B1(G559), .B2(new_n551), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT83), .ZN(G148));
  NAND2_X1  g188(.A1(new_n550), .A2(new_n606), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n602), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g192(.A(new_n468), .B1(new_n458), .B2(new_n459), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n479), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n481), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n623), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n633), .B2(new_n634), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n636), .B(new_n640), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT86), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n622), .ZN(new_n655));
  NOR2_X1   g230(.A1(G2072), .A2(G2078), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n442), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n678), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  NAND2_X1  g256(.A1(new_n479), .A2(G141), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n481), .A2(G129), .ZN(new_n683));
  NAND3_X1  g258(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT26), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  AOI22_X1  g262(.A1(G105), .A2(new_n468), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(G32), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT27), .B(G1996), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G5), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G171), .B2(new_n696), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(G1961), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G164), .A2(new_n691), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G27), .B2(new_n691), .ZN(new_n701));
  INV_X1    g276(.A(G2078), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n698), .A2(G1961), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n693), .B2(new_n694), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n699), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT31), .B(G11), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n628), .A2(new_n691), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT97), .B(G28), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(KEYINPUT30), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n709), .B2(KEYINPUT30), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n707), .B(new_n708), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n691), .A2(G33), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n479), .A2(G139), .ZN(new_n714));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n715));
  INV_X1    g290(.A(G127), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n460), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2105), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n714), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n713), .B1(new_n722), .B2(new_n691), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT24), .B(G34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(new_n691), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT95), .Z(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n477), .B2(new_n691), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n723), .A2(G2072), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n712), .B(new_n729), .C1(G2072), .C2(new_n723), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n724), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT96), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n696), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n696), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1966), .ZN(new_n735));
  NOR4_X1   g310(.A1(new_n706), .A2(new_n730), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n691), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n481), .A2(G128), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n475), .A2(G116), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n479), .A2(G140), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n740), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n740), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n738), .B1(new_n749), .B2(new_n691), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2067), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n691), .A2(G35), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT98), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n691), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G2090), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT100), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G4), .A2(G16), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n603), .B2(G16), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G1348), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(G1348), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT89), .B(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G20), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT101), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G16), .B2(G299), .ZN(new_n768));
  INV_X1    g343(.A(G1956), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n762), .A2(new_n763), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n701), .A2(new_n702), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n764), .A2(G19), .ZN(new_n773));
  INV_X1    g348(.A(new_n550), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n764), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n756), .A2(G2090), .B1(new_n775), .B2(G1341), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n772), .B(new_n776), .C1(G1341), .C2(new_n775), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n736), .A2(new_n759), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  MUX2_X1   g353(.A(G303), .B(G22), .S(new_n764), .Z(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n696), .A2(G6), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G305), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT32), .B(G1981), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT91), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n785), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n781), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n696), .A2(G23), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n696), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT33), .B(G1976), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT92), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n788), .A2(KEYINPUT34), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT34), .B1(new_n788), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n479), .A2(G131), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n481), .A2(G119), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n475), .A2(G107), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G25), .B(new_n801), .S(G29), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT88), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G290), .B(G24), .S(new_n764), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT90), .B(G1986), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n795), .A2(new_n796), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT36), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(KEYINPUT36), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n778), .B1(new_n812), .B2(new_n813), .ZN(G311));
  XNOR2_X1  g389(.A(G311), .B(KEYINPUT102), .ZN(G150));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n531), .A2(new_n816), .B1(new_n526), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT103), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(new_n509), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(KEYINPUT104), .A3(new_n821), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n774), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n823), .A3(new_n550), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n603), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n822), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  OAI21_X1  g412(.A(new_n689), .B1(new_n747), .B2(new_n748), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n740), .A2(new_n745), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT94), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n840), .A2(new_n690), .A3(new_n746), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n487), .B1(new_n474), .B2(new_n490), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n494), .B(new_n497), .C1(new_n842), .C2(new_n489), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n838), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n838), .B2(new_n841), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n721), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n843), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n747), .A2(new_n748), .A3(new_n689), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n690), .B1(new_n840), .B2(new_n746), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n838), .A2(new_n841), .A3(new_n843), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n722), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n801), .B(new_n620), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n481), .A2(G130), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G142), .B2(new_n479), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n854), .B(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n846), .A2(new_n852), .A3(new_n853), .A4(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(new_n485), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT105), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n628), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n846), .B2(new_n852), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n853), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n846), .A2(new_n852), .A3(new_n860), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n864), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n867), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT107), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n869), .A2(new_n864), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n846), .A2(new_n852), .ZN(new_n876));
  INV_X1    g451(.A(new_n860), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(KEYINPUT106), .A3(new_n869), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n861), .A2(new_n865), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n874), .A2(new_n884), .A3(KEYINPUT40), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT40), .B1(new_n874), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(G395));
  XNOR2_X1  g462(.A(new_n828), .B(new_n615), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n602), .A2(G299), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n602), .A2(G299), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n893));
  INV_X1    g468(.A(new_n891), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n889), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT41), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G305), .B(G303), .ZN(new_n899));
  XNOR2_X1  g474(.A(G290), .B(KEYINPUT109), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G288), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n790), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n899), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n904), .A3(new_n899), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n898), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n822), .A2(new_n606), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  XNOR2_X1  g490(.A(G168), .B(G301), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n826), .A2(new_n827), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n826), .B2(new_n827), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n895), .A2(new_n896), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n890), .A2(new_n891), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n908), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n871), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n906), .A2(KEYINPUT110), .A3(new_n907), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  INV_X1    g502(.A(new_n907), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n905), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n920), .B2(new_n923), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n893), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n894), .A2(new_n889), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n922), .B2(KEYINPUT41), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n918), .A2(new_n919), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n923), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n926), .A3(new_n929), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n871), .A4(new_n924), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n925), .B2(new_n931), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n871), .A3(new_n924), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n939), .ZN(new_n944));
  MUX2_X1   g519(.A(new_n941), .B(new_n944), .S(KEYINPUT44), .Z(G397));
  XOR2_X1   g520(.A(KEYINPUT111), .B(G1384), .Z(new_n946));
  NAND2_X1  g521(.A1(new_n843), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n469), .A2(new_n950), .A3(G40), .A4(new_n476), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n472), .A2(new_n463), .ZN(new_n952));
  NAND2_X1  g527(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n461), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n462), .A2(new_n463), .ZN(new_n955));
  OAI21_X1  g530(.A(G2105), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n468), .A2(G101), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n476), .A2(new_n956), .A3(G40), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT113), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n749), .B(G2067), .ZN(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n689), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n801), .A2(new_n805), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n801), .A2(new_n805), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(G1986), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(G1341), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n494), .A2(new_n497), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n492), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n843), .A2(KEYINPUT114), .A3(new_n973), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n960), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT45), .B(new_n946), .C1(new_n492), .C2(new_n974), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(new_n959), .A3(new_n951), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n500), .A2(new_n973), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(new_n948), .ZN(new_n985));
  AOI22_X1  g560(.A1(KEYINPUT124), .A2(new_n981), .B1(new_n985), .B2(new_n963), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT124), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n960), .B1(new_n978), .B2(new_n977), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(new_n972), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT125), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n979), .A2(new_n980), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(KEYINPUT124), .A3(new_n971), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n984), .A2(new_n948), .ZN(new_n993));
  INV_X1    g568(.A(new_n983), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(new_n963), .ZN(new_n995));
  AND4_X1   g570(.A1(KEYINPUT125), .A2(new_n992), .A3(new_n989), .A4(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n774), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n977), .A2(KEYINPUT50), .A3(new_n978), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n980), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n500), .A2(new_n1003), .A3(new_n973), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n1000), .B2(new_n980), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n769), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G299), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n564), .A2(G91), .B1(G651), .B2(new_n568), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(new_n1009), .A3(new_n1010), .A4(new_n560), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n985), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT61), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1007), .A2(new_n1017), .A3(KEYINPUT61), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n978), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT114), .B1(new_n843), .B2(new_n973), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1003), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n980), .ZN(new_n1027));
  INV_X1    g602(.A(G1348), .ZN(new_n1028));
  INV_X1    g603(.A(G2067), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1027), .A2(new_n1028), .B1(new_n1029), .B2(new_n988), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT60), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n602), .B1(new_n1030), .B2(KEYINPUT60), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT59), .B(new_n774), .C1(new_n990), .C2(new_n996), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n999), .A2(new_n1022), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT126), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n1038));
  OR3_X1    g613(.A1(new_n1030), .A2(new_n1038), .A3(new_n602), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1030), .B2(new_n602), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n985), .A2(new_n1016), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1007), .A2(new_n1042), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1018), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1036), .A2(new_n1037), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n790), .A2(G1976), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n991), .A2(new_n1047), .A3(new_n1049), .A4(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT117), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n988), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n586), .A2(new_n1056), .A3(new_n587), .ZN(new_n1057));
  INV_X1    g632(.A(G86), .ZN(new_n1058));
  OAI221_X1 g633(.A(new_n582), .B1(new_n1058), .B2(new_n526), .C1(new_n584), .C2(new_n509), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT49), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1051), .A2(new_n1055), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n991), .A2(new_n1047), .A3(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT116), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1067), .A3(KEYINPUT52), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n960), .B1(new_n979), .B2(new_n1003), .ZN(new_n1070));
  INV_X1    g645(.A(G2090), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1026), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n993), .A2(new_n994), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n780), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(G166), .B2(new_n1052), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1076), .A2(KEYINPUT115), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT115), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1081), .A3(G8), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1063), .A2(new_n1069), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1005), .A2(G2090), .A3(new_n1006), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1074), .ZN(new_n1087));
  OAI21_X1  g662(.A(G8), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT53), .B1(new_n985), .B2(new_n702), .ZN(new_n1090));
  INV_X1    g665(.A(G1961), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1091), .B2(new_n1027), .ZN(new_n1092));
  INV_X1    g667(.A(new_n948), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n500), .A2(new_n973), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n980), .B(new_n1094), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n702), .A2(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(G171), .B(KEYINPUT54), .Z(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT53), .B1(KEYINPUT127), .B2(G2078), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1099), .B(new_n958), .C1(KEYINPUT127), .C2(G2078), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1100), .A2(new_n982), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n949), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1097), .A2(new_n1098), .B1(new_n1092), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  INV_X1    g679(.A(G1966), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1095), .A2(KEYINPUT119), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1070), .A2(new_n724), .A3(new_n1026), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT119), .B1(new_n1095), .B2(new_n1105), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1052), .B1(new_n1110), .B2(G168), .ZN(new_n1111));
  OAI21_X1  g686(.A(G286), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1104), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1109), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(G168), .A3(new_n1107), .A4(new_n1106), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1115), .A2(new_n1104), .A3(G8), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1089), .B(new_n1103), .C1(new_n1113), .C2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1045), .A2(new_n1046), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT62), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1063), .A2(new_n1069), .A3(new_n1082), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1088), .A2(new_n1078), .A3(new_n1076), .ZN(new_n1121));
  AND4_X1   g696(.A1(G171), .A2(new_n1120), .A3(new_n1121), .A4(new_n1097), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1116), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(new_n1115), .A3(G8), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT51), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(G1976), .B(G288), .C1(new_n1062), .C2(new_n1053), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1057), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1053), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1082), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1110), .A2(new_n1052), .A3(G286), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1120), .A2(new_n1134), .A3(new_n1121), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1075), .A2(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1085), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1120), .A2(new_n1134), .A3(KEYINPUT63), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n969), .B1(new_n1118), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n749), .A2(new_n1029), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n962), .A2(new_n964), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n966), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1146), .A2(new_n961), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n961), .A2(new_n963), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT46), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n962), .A2(new_n690), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n961), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT47), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n967), .A2(new_n961), .ZN(new_n1153));
  NOR4_X1   g728(.A1(G290), .A2(new_n949), .A3(new_n960), .A4(G1986), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT48), .Z(new_n1155));
  AOI211_X1 g730(.A(new_n1147), .B(new_n1152), .C1(new_n1153), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g732(.A1(new_n874), .A2(new_n884), .ZN(new_n1159));
  INV_X1    g733(.A(G227), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n645), .A2(new_n1160), .A3(G319), .ZN(new_n1161));
  AOI21_X1  g735(.A(new_n1161), .B1(new_n679), .B2(new_n680), .ZN(new_n1162));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n941), .A3(new_n1162), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


