//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT65), .A3(G137), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT65), .B1(new_n187), .B2(G137), .ZN(new_n192));
  OAI21_X1  g006(.A(G131), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n187), .A2(G137), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(G134), .B2(new_n189), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n187), .A2(KEYINPUT11), .A3(G137), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n194), .B(new_n195), .C1(new_n197), .C2(new_n198), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n193), .A2(new_n199), .A3(KEYINPUT66), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n193), .B2(new_n199), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT64), .A3(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G128), .ZN(new_n214));
  AOI221_X4 g028(.A(new_n202), .B1(new_n203), .B2(new_n205), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n214), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n205), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT67), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n200), .A2(new_n201), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n203), .A2(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G131), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n199), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT2), .B(G113), .Z(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n219), .A2(KEYINPUT70), .A3(new_n230), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n231), .A2(new_n240), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n219), .A2(new_n241), .A3(new_n230), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT28), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  INV_X1    g067(.A(G237), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n253), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(G902), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n216), .A2(new_n217), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n199), .A3(new_n193), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n230), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n240), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n244), .B1(new_n247), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n243), .B2(new_n244), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n267), .A2(new_n268), .A3(new_n257), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n267), .B2(new_n257), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n247), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT30), .B1(new_n230), .B2(new_n263), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n241), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n226), .B2(new_n229), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n219), .A2(KEYINPUT68), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT68), .B1(new_n219), .B2(new_n276), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT69), .B(new_n274), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n272), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n259), .B1(new_n283), .B2(new_n257), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n261), .B1(new_n271), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G472), .ZN(new_n286));
  INV_X1    g100(.A(new_n267), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n258), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n282), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n247), .A2(new_n257), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT31), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n293), .B(new_n290), .C1(new_n281), .C2(new_n282), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n288), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n219), .A2(new_n276), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n219), .A2(KEYINPUT68), .A3(new_n276), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT69), .B1(new_n306), .B2(new_n274), .ZN(new_n307));
  INV_X1    g121(.A(new_n282), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n291), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n293), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n290), .B1(new_n281), .B2(new_n282), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT31), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n310), .A2(new_n312), .B1(new_n287), .B2(new_n258), .ZN(new_n313));
  INV_X1    g127(.A(new_n297), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT32), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n286), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n301), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  OR3_X1    g138(.A1(new_n322), .A2(new_n324), .A3(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(G146), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n323), .B2(new_n325), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n210), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n234), .B2(G128), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n337), .B(new_n338), .C1(G119), .C2(new_n204), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G110), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT73), .Z(new_n341));
  XOR2_X1   g155(.A(KEYINPUT24), .B(G110), .Z(new_n342));
  XNOR2_X1  g156(.A(G119), .B(G128), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n327), .A2(KEYINPUT75), .A3(G146), .A4(new_n329), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n335), .A2(new_n341), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n339), .A2(G110), .B1(new_n343), .B2(new_n342), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n321), .A2(new_n210), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n330), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT76), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n355), .B(KEYINPUT22), .Z(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n189), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n351), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n350), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n363));
  INV_X1    g177(.A(G217), .ZN(new_n364));
  INV_X1    g178(.A(G902), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(G234), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n360), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n366), .A2(G902), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT79), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n320), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n254), .A2(new_n255), .A3(G214), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(G143), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT93), .B1(new_n378), .B2(new_n194), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(new_n207), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G131), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n379), .A2(new_n382), .B1(new_n194), .B2(new_n378), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n335), .A2(new_n345), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(KEYINPUT17), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n388));
  OAI211_X1 g202(.A(KEYINPUT18), .B(G131), .C1(new_n380), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n388), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n348), .B1(new_n326), .B2(new_n210), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n380), .A2(new_n388), .A3(KEYINPUT18), .A4(G131), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G113), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(G104), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT95), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n387), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n394), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n385), .B2(new_n386), .ZN(new_n400));
  INV_X1    g214(.A(new_n396), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n365), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT96), .B(G475), .Z(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT19), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n321), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n326), .B2(new_n407), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n330), .B1(G146), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n394), .B1(new_n410), .B2(new_n383), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n396), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT94), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n414), .A3(new_n396), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n413), .A2(new_n415), .B1(new_n400), .B2(new_n397), .ZN(new_n416));
  NOR2_X1   g230(.A1(G475), .A2(G902), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n416), .A2(KEYINPUT20), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n415), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n414), .B1(new_n411), .B2(new_n396), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n398), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n406), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT97), .B1(new_n204), .B2(G143), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n207), .A3(G128), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n427), .A2(new_n429), .B1(new_n204), .B2(G143), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n187), .ZN(new_n431));
  INV_X1    g245(.A(G122), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G116), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(G116), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G107), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(KEYINPUT98), .A3(KEYINPUT14), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT14), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT98), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n433), .B2(new_n440), .ZN(new_n443));
  AND4_X1   g257(.A1(new_n435), .A2(new_n439), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n431), .B(new_n438), .C1(new_n444), .C2(new_n437), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n436), .B(new_n437), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT13), .B1(new_n204), .B2(G143), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n187), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n430), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT9), .B(G234), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n453), .A2(new_n364), .A3(G953), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n450), .A3(new_n454), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT99), .A3(new_n457), .ZN(new_n458));
  OR3_X1    g272(.A1(new_n451), .A2(KEYINPUT99), .A3(new_n455), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT100), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n461), .A3(new_n365), .A4(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n459), .A3(new_n365), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n466), .B2(KEYINPUT100), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(KEYINPUT100), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT101), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT101), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n465), .B(new_n471), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n426), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G952), .ZN(new_n474));
  AOI211_X1 g288(.A(G953), .B(new_n474), .C1(G234), .C2(G237), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT21), .B(G898), .Z(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n365), .B(new_n255), .C1(G234), .C2(G237), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n225), .A2(G125), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(G125), .B2(new_n262), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G224), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(G953), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n490), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n492), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n495));
  XOR2_X1   g309(.A(G110), .B(G122), .Z(new_n496));
  INV_X1    g310(.A(G104), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT3), .B1(new_n497), .B2(G107), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n437), .A3(G104), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(G107), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(G101), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n502), .A2(new_n506), .A3(new_n503), .A4(G101), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n503), .B1(new_n502), .B2(G101), .ZN(new_n509));
  INV_X1    g323(.A(G101), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n498), .A2(new_n500), .A3(new_n510), .A4(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n240), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n514));
  INV_X1    g328(.A(new_n501), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n497), .A2(G107), .ZN(new_n516));
  OAI21_X1  g330(.A(G101), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n511), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n238), .A2(new_n239), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT5), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(G113), .C1(KEYINPUT5), .C2(new_n235), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n513), .A2(new_n514), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n514), .B1(new_n513), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n496), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n496), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n513), .A2(new_n527), .A3(new_n523), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n495), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n513), .A2(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT87), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n513), .A2(new_n514), .A3(new_n523), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT6), .B1(new_n533), .B2(new_n496), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n494), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G210), .B1(G237), .B2(G902), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT7), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n528), .B1(new_n493), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n522), .A2(new_n520), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT90), .B1(new_n539), .B2(new_n518), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(new_n523), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n523), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT89), .B(KEYINPUT8), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n496), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n484), .B1(new_n537), .B2(new_n490), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n365), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n535), .A2(new_n536), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n536), .B1(new_n535), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n482), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G140), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n255), .A2(G227), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n215), .A2(new_n218), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT83), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT10), .A4(new_n519), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n505), .A2(new_n507), .B1(new_n511), .B2(new_n509), .ZN(new_n559));
  MUX2_X1   g373(.A(new_n214), .B(new_n205), .S(new_n203), .Z(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n519), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n559), .A2(new_n226), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT10), .B(new_n519), .C1(new_n215), .C2(new_n218), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT83), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n229), .ZN(new_n567));
  INV_X1    g381(.A(new_n229), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n558), .A2(new_n568), .A3(new_n563), .A4(new_n565), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n555), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n555), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n518), .A2(new_n216), .A3(new_n217), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n568), .B1(new_n561), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT12), .B1(new_n229), .B2(KEYINPUT84), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n578));
  INV_X1    g392(.A(G469), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n577), .A2(new_n365), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n571), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT85), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n571), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n567), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n575), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n569), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n555), .B(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n583), .B1(new_n593), .B2(new_n579), .ZN(new_n594));
  OAI21_X1  g408(.A(G221), .B1(new_n453), .B2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n481), .A2(new_n552), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n376), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n295), .A2(new_n297), .ZN(new_n600));
  OAI21_X1  g414(.A(G472), .B1(new_n313), .B2(G902), .ZN(new_n601));
  AND4_X1   g415(.A1(new_n600), .A2(new_n601), .A3(new_n595), .A4(new_n594), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n375), .A2(new_n479), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n552), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n458), .A2(new_n459), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n457), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n457), .A2(new_n609), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(KEYINPUT33), .A3(new_n456), .A4(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n608), .A2(new_n612), .A3(G478), .A4(new_n365), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n466), .A2(new_n462), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n426), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n536), .ZN(new_n617));
  INV_X1    g431(.A(new_n494), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n619));
  INV_X1    g433(.A(new_n528), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT6), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n526), .A2(new_n495), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n617), .B1(new_n623), .B2(new_n548), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n535), .A2(new_n536), .A3(new_n549), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(KEYINPUT102), .A3(new_n482), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n606), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G6));
  AOI21_X1  g446(.A(new_n404), .B1(new_n402), .B2(new_n365), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n420), .B1(new_n416), .B2(new_n418), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n424), .A2(new_n421), .A3(new_n417), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n470), .A2(new_n636), .A3(new_n472), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n606), .A3(new_n627), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n604), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT35), .B(G107), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NOR2_X1   g455(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n350), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n373), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n370), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n597), .A2(new_n600), .A3(new_n601), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT37), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(G110), .Z(G12));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n475), .B1(new_n478), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n594), .A2(new_n595), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n638), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n653), .A2(new_n301), .A3(new_n319), .A4(new_n645), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n318), .B1(new_n317), .B2(new_n286), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(KEYINPUT105), .A3(new_n645), .A4(new_n653), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  INV_X1    g476(.A(KEYINPUT38), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n626), .B(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n370), .A2(new_n644), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n482), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n426), .A2(new_n470), .A3(new_n472), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n665), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n666), .A2(KEYINPUT107), .A3(new_n668), .A4(new_n482), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n664), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n650), .B(KEYINPUT39), .ZN(new_n673));
  OR3_X1    g487(.A1(new_n596), .A2(KEYINPUT108), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT108), .B1(new_n596), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n248), .A2(new_n258), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT106), .Z(new_n680));
  OAI21_X1  g494(.A(new_n365), .B1(new_n680), .B2(new_n311), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n317), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n674), .A2(KEYINPUT40), .A3(new_n675), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n672), .A2(new_n678), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n628), .A2(new_n652), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n659), .A2(new_n687), .A3(new_n645), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(new_n301), .A3(new_n319), .A4(new_n645), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  AND2_X1   g507(.A1(new_n370), .A2(new_n374), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n626), .B2(new_n482), .ZN(new_n695));
  INV_X1    g509(.A(new_n482), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n605), .B(new_n696), .C1(new_n624), .C2(new_n625), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n426), .A2(new_n615), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n694), .A2(new_n301), .A3(new_n319), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n365), .B1(new_n570), .B2(new_n576), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n583), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n595), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n479), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT41), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G113), .ZN(G15));
  NAND4_X1  g522(.A1(new_n301), .A2(new_n319), .A3(new_n694), .A4(new_n705), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(new_n638), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NOR2_X1   g525(.A1(new_n703), .A2(new_n704), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n606), .A3(new_n627), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n301), .A2(new_n713), .A3(new_n319), .A4(new_n645), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(new_n481), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  OAI22_X1  g530(.A1(new_n292), .A2(new_n294), .B1(new_n257), .B2(new_n251), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n297), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n694), .A2(new_n705), .A3(new_n601), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n668), .A2(new_n606), .A3(new_n627), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n695), .A2(new_n697), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(KEYINPUT110), .A3(new_n668), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n719), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n432), .ZN(G24));
  AND2_X1   g540(.A1(new_n601), .A2(new_n718), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n616), .ZN(new_n728));
  INV_X1    g542(.A(new_n723), .ZN(new_n729));
  INV_X1    g543(.A(new_n712), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n645), .A2(new_n651), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n324), .ZN(G27));
  INV_X1    g547(.A(new_n626), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n482), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n596), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n320), .A2(new_n375), .A3(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n698), .A2(KEYINPUT42), .A3(new_n650), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n375), .B1(new_n317), .B2(new_n286), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n698), .A2(new_n650), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n736), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n738), .A2(new_n739), .B1(KEYINPUT42), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  AND2_X1   g558(.A1(new_n637), .A2(new_n651), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n588), .A2(new_n592), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n588), .A2(KEYINPUT45), .A3(new_n592), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(G469), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n579), .A2(new_n365), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n748), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n753), .B(KEYINPUT46), .C1(new_n579), .C2(new_n365), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n583), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n673), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n595), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT111), .Z(new_n761));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n666), .B1(new_n600), .B2(new_n601), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n406), .B(new_n615), .C1(new_n419), .C2(new_n425), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT20), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n424), .A2(new_n765), .A3(new_n417), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n633), .B1(new_n634), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT43), .B1(new_n767), .B2(KEYINPUT112), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n426), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n764), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT113), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n771), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n762), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n735), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n763), .A2(new_n777), .A3(KEYINPUT114), .A4(KEYINPUT44), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT115), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n779), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n786), .A3(new_n781), .A4(new_n782), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n761), .A2(new_n784), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND2_X1  g603(.A1(new_n758), .A2(new_n595), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n659), .A2(new_n735), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n375), .A3(new_n741), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NOR2_X1   g609(.A1(G952), .A2(G953), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT121), .ZN(new_n797));
  INV_X1    g611(.A(new_n683), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n730), .A2(new_n735), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n694), .A3(new_n799), .A4(new_n475), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n426), .A3(new_n615), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n694), .A2(new_n777), .A3(new_n475), .A4(new_n727), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n712), .ZN(new_n804));
  INV_X1    g618(.A(new_n664), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n482), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n802), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(KEYINPUT50), .A3(new_n712), .A4(new_n806), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n801), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n703), .B(KEYINPUT116), .Z(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT120), .Z(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n595), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n781), .B(new_n803), .C1(new_n792), .C2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n777), .A2(new_n475), .A3(new_n799), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n645), .A3(new_n727), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n810), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n255), .A2(G952), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n815), .A2(new_n740), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT48), .Z(new_n823));
  NOR4_X1   g637(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n800), .A2(new_n698), .ZN(new_n825));
  INV_X1    g639(.A(new_n732), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n798), .A2(new_n652), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n722), .A2(new_n724), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n666), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n661), .A2(new_n692), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n732), .B1(new_n656), .B2(new_n660), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .A3(new_n692), .A4(new_n829), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n604), .ZN(new_n836));
  INV_X1    g650(.A(new_n469), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n698), .B1(new_n426), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n836), .A2(new_n482), .A3(new_n626), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n598), .A2(new_n839), .A3(new_n646), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n725), .B1(new_n700), .B2(new_n705), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT117), .A3(new_n710), .A4(new_n715), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n481), .A2(new_n714), .B1(new_n709), .B2(new_n638), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n694), .A2(new_n705), .A3(new_n601), .A4(new_n718), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT110), .B1(new_n723), .B2(new_n668), .ZN(new_n846));
  AND4_X1   g660(.A1(KEYINPUT110), .A2(new_n668), .A3(new_n606), .A4(new_n627), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n705), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n301), .A2(new_n319), .A3(new_n694), .A4(new_n699), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n843), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n840), .B1(new_n842), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n301), .A2(new_n319), .A3(new_n837), .A4(new_n636), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n728), .ZN(new_n856));
  INV_X1    g670(.A(new_n731), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n736), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n738), .A2(new_n739), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n854), .A2(new_n858), .A3(new_n859), .A4(new_n746), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT53), .B1(new_n835), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n842), .A2(new_n852), .ZN(new_n863));
  INV_X1    g677(.A(new_n840), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n832), .A2(new_n866), .A3(new_n834), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n833), .A2(new_n692), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT118), .A3(KEYINPUT52), .A4(new_n829), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n865), .A2(new_n867), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n871), .A3(KEYINPUT54), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n868), .B1(new_n835), .B2(new_n861), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n743), .A2(KEYINPUT53), .A3(new_n746), .A4(new_n858), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n841), .A2(new_n710), .A3(new_n715), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n840), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n867), .A2(new_n870), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n824), .A2(new_n825), .A3(new_n872), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n804), .A2(new_n729), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n797), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n694), .A2(new_n482), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n774), .B1(new_n811), .B2(KEYINPUT49), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(KEYINPUT49), .B2(new_n811), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n805), .A2(new_n704), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n798), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n884), .B2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n255), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n365), .B1(new_n873), .B2(new_n877), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n529), .A2(new_n534), .A3(new_n494), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n623), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n891), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n867), .A2(new_n870), .A3(new_n876), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n832), .A2(new_n834), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n865), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(G902), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n873), .A2(new_n877), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT122), .A3(G902), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n617), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n897), .B1(new_n906), .B2(new_n908), .ZN(G51));
  OAI21_X1  g723(.A(new_n878), .B1(new_n898), .B2(new_n900), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n880), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n755), .B(KEYINPUT123), .Z(new_n912));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n577), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n903), .A2(new_n754), .A3(new_n905), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n890), .B1(new_n917), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n903), .A2(new_n905), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n416), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n903), .A2(new_n905), .A3(new_n424), .A4(new_n920), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n891), .A3(new_n923), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n910), .B2(new_n880), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n608), .A2(new_n612), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n927), .A2(KEYINPUT124), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT124), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n872), .B2(new_n880), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n891), .B1(new_n931), .B2(new_n928), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(G63));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n904), .A2(new_n643), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n891), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n873), .B2(new_n877), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n371), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n934), .B(KEYINPUT61), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n941), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n890), .B1(new_n940), .B2(new_n643), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n942), .A2(new_n947), .ZN(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n477), .B2(new_n489), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n853), .B2(G953), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n621), .B(new_n622), .C1(G898), .C2(new_n255), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  INV_X1    g766(.A(new_n306), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(new_n273), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n409), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n794), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n869), .A2(KEYINPUT62), .A3(new_n685), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n833), .A2(new_n692), .ZN(new_n960));
  INV_X1    g774(.A(new_n685), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n596), .A2(new_n673), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n376), .A2(new_n964), .A3(new_n781), .A4(new_n838), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n788), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(KEYINPUT126), .B(new_n956), .C1(new_n967), .C2(G953), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  AOI21_X1  g783(.A(G953), .B1(new_n963), .B2(new_n966), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n955), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n761), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n828), .A2(new_n740), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n869), .A2(new_n794), .A3(new_n743), .A4(new_n746), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n255), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(G900), .B2(new_n255), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n979), .B(new_n982), .C1(G900), .C2(new_n255), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n955), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n972), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n973), .B1(new_n972), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(new_n283), .A2(new_n258), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n977), .A2(new_n978), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n853), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n890), .ZN(new_n994));
  INV_X1    g808(.A(new_n992), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n283), .A2(new_n258), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n862), .A2(new_n871), .A3(new_n997), .A4(new_n988), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n995), .B1(new_n967), .B2(new_n853), .ZN(new_n999));
  OAI221_X1 g813(.A(new_n994), .B1(new_n995), .B2(new_n998), .C1(new_n999), .C2(new_n997), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(G57));
endmodule


