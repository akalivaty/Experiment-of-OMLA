//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(KEYINPUT66), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(KEYINPUT66), .B2(new_n457), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n461), .A2(new_n463), .A3(new_n467), .A4(G125), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n460), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n461), .ZN(new_n474));
  NOR3_X1   g049(.A1(new_n473), .A2(G2105), .A3(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n469), .A2(G2105), .B1(new_n475), .B2(G137), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND4_X1   g055(.A1(new_n477), .A2(new_n470), .A3(new_n472), .A4(new_n479), .ZN(new_n481));
  OAI21_X1  g056(.A(G101), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(KEYINPUT70), .B(G101), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n476), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  NAND2_X1  g063(.A1(new_n470), .A2(new_n472), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n474), .B1(new_n489), .B2(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G124), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT72), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT73), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n475), .A2(G136), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n473), .A2(new_n479), .A3(new_n474), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(new_n499), .A3(G124), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n493), .A2(new_n496), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  AND3_X1   g077(.A1(new_n479), .A2(G102), .A3(G2104), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n479), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n490), .A2(KEYINPUT4), .A3(G138), .A4(new_n479), .ZN(new_n507));
  NAND2_X1  g082(.A1(G114), .A2(G2104), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n490), .B2(G126), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n506), .B(new_n507), .C1(new_n510), .C2(new_n479), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n520), .A2(G651), .B1(new_n524), .B2(G50), .ZN(new_n525));
  OR3_X1    g100(.A1(new_n518), .A2(new_n523), .A3(KEYINPUT74), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n518), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n524), .A2(G51), .ZN(new_n532));
  INV_X1    g107(.A(new_n528), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n515), .A2(new_n517), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT75), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  AND4_X1   g114(.A1(new_n532), .A2(new_n534), .A3(new_n537), .A4(new_n539), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n518), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n524), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n533), .A2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n518), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(new_n524), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  AOI22_X1  g136(.A1(new_n535), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G651), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n526), .A2(G91), .A3(new_n527), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(new_n524), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n564), .A2(new_n565), .A3(new_n569), .A4(new_n570), .ZN(G299));
  NAND4_X1  g146(.A1(new_n534), .A2(new_n532), .A3(new_n537), .A4(new_n539), .ZN(G286));
  NAND3_X1  g147(.A1(new_n526), .A2(G87), .A3(new_n527), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n524), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n524), .A2(G48), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n535), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n563), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT77), .B1(new_n528), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n526), .A2(new_n582), .A3(G86), .A4(new_n527), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n533), .A2(G85), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT78), .B(G47), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n563), .B2(new_n587), .C1(new_n567), .C2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n528), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n518), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n524), .B2(G54), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT10), .B1(new_n528), .B2(new_n591), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G321));
  MUX2_X1   g176(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g178(.A(KEYINPUT79), .B(G559), .Z(new_n604));
  OAI21_X1  g179(.A(new_n599), .B1(G860), .B2(new_n604), .ZN(G148));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g184(.A1(new_n480), .A2(new_n481), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n610), .A2(new_n461), .A3(new_n463), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT80), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n498), .A2(G123), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n475), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n479), .B2(G111), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n633), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n631), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n637), .A2(new_n640), .A3(new_n642), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT82), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n644), .A2(new_n648), .A3(G14), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  AOI21_X1  g236(.A(KEYINPUT18), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n674), .C2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT84), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n681), .B(new_n684), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G35), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G162), .B2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT97), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(KEYINPUT97), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(G2090), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G19), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n555), .B2(new_n698), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(G1341), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(G1341), .ZN(new_n702));
  OR2_X1    g277(.A1(G5), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G301), .B2(new_n698), .ZN(new_n704));
  INV_X1    g279(.A(G1961), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n701), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(G299), .A2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n698), .A2(G20), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1956), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G32), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n610), .A2(G105), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n475), .A2(G141), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n498), .A2(G129), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n707), .A2(new_n714), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n695), .B2(new_n696), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n479), .ZN(new_n731));
  INV_X1    g306(.A(G139), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT91), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n461), .A2(new_n463), .A3(G127), .ZN(new_n735));
  INV_X1    g310(.A(G115), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n462), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2105), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n687), .A2(G33), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(KEYINPUT92), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n743), .A2(G2072), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n743), .A2(new_n745), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(G2072), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n697), .A2(new_n728), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n624), .A2(KEYINPUT95), .A3(G29), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n622), .A2(new_n623), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n687), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G28), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n687), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n698), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1966), .Z(new_n764));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n704), .A2(new_n705), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n761), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n755), .A2(new_n766), .A3(new_n756), .A4(new_n760), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n763), .B(G1966), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT96), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n691), .A2(G2090), .A3(new_n694), .ZN(new_n772));
  AND2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  NOR2_X1   g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n687), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(KEYINPUT93), .B2(G2084), .C1(new_n487), .C2(new_n687), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT93), .A2(G2084), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n776), .B(new_n777), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n498), .A2(G128), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n475), .A2(G140), .ZN(new_n780));
  NOR2_X1   g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(new_n479), .B2(G116), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n687), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n771), .A2(new_n772), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n750), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n698), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n698), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G1971), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n698), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n698), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT33), .B(G1976), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT88), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n801), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n794), .A2(G1971), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n795), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n698), .A2(G6), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n584), .B2(new_n698), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(new_n683), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n683), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n805), .B(new_n812), .C1(new_n809), .C2(new_n810), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(KEYINPUT89), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n687), .A2(G25), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n498), .A2(G119), .ZN(new_n820));
  OR2_X1    g395(.A1(G95), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n822));
  INV_X1    g397(.A(G131), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n820), .B(new_n822), .C1(new_n823), .C2(new_n731), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(new_n687), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT85), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT35), .B(G1991), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n698), .A2(G24), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G290), .B2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT86), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(G1986), .Z(new_n833));
  NAND4_X1  g408(.A1(new_n816), .A2(new_n818), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(new_n814), .A3(new_n815), .A4(new_n829), .ZN(new_n835));
  INV_X1    g410(.A(new_n818), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n817), .A2(KEYINPUT89), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n792), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G4), .A2(G16), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n599), .B2(G16), .ZN(new_n841));
  INV_X1    g416(.A(G1348), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n687), .A2(G27), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G164), .B2(new_n687), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G2078), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n839), .A2(KEYINPUT100), .A3(new_n843), .A4(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n792), .A2(new_n834), .A3(new_n838), .A4(new_n843), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(G311));
  NAND3_X1  g427(.A1(new_n839), .A2(new_n843), .A3(new_n847), .ZN(G150));
  AOI22_X1  g428(.A1(new_n535), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n563), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n524), .A2(G55), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n855), .B(new_n856), .C1(new_n528), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n599), .A2(G559), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT38), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT39), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(KEYINPUT101), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n554), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n555), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n863), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n860), .B1(new_n870), .B2(G860), .ZN(G145));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n734), .A2(new_n722), .A3(new_n738), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n722), .B1(new_n738), .B2(new_n734), .ZN(new_n875));
  XNOR2_X1  g450(.A(G164), .B(new_n783), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n498), .A2(G130), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n475), .A2(G142), .ZN(new_n882));
  NOR2_X1   g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(new_n479), .B2(G118), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n613), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n613), .A2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n824), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n613), .A2(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n825), .A3(new_n886), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n877), .A2(new_n893), .A3(new_n878), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n880), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n753), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n753), .A2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n487), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n624), .A2(KEYINPUT102), .ZN(new_n901));
  NAND3_X1  g476(.A1(G160), .A2(new_n901), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n501), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n902), .A3(G162), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n895), .B(new_n906), .C1(new_n880), .C2(new_n892), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n879), .A2(new_n892), .A3(KEYINPUT104), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT104), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n877), .A3(new_n878), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n908), .A2(new_n905), .A3(new_n904), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n872), .B(new_n907), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g491(.A1(new_n858), .A2(G868), .ZN(new_n917));
  XNOR2_X1  g492(.A(G288), .B(G303), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G290), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n584), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT42), .Z(new_n921));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n869), .B(new_n606), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n598), .B(G299), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT41), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n923), .A2(new_n924), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n929), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n921), .B(new_n922), .C1(new_n933), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n917), .B1(new_n935), .B2(G868), .ZN(G295));
  AOI21_X1  g511(.A(new_n917), .B1(new_n935), .B2(G868), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g513(.A1(G286), .A2(KEYINPUT107), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(G286), .A2(KEYINPUT107), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(G171), .ZN(new_n942));
  OR2_X1    g517(.A1(G286), .A2(KEYINPUT107), .ZN(new_n943));
  AOI21_X1  g518(.A(G301), .B1(new_n943), .B2(new_n939), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n869), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(G171), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(G301), .A3(new_n939), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n868), .A4(new_n865), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n927), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n928), .A2(new_n948), .A3(new_n945), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n938), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n928), .A2(new_n948), .A3(new_n945), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n920), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n920), .B1(new_n953), .B2(new_n955), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT43), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n927), .B1(new_n945), .B2(new_n948), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT108), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n962), .B(new_n957), .C1(KEYINPUT108), .C2(new_n954), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n920), .B1(new_n954), .B2(new_n961), .ZN(new_n964));
  AND4_X1   g539(.A1(KEYINPUT43), .A2(new_n963), .A3(new_n872), .A4(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n958), .B2(new_n959), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n968), .A2(new_n963), .A3(new_n872), .A4(new_n964), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT4), .B(new_n461), .C1(new_n478), .C2(new_n460), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n479), .A2(G138), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n506), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(G126), .B(new_n461), .C1(new_n478), .C2(new_n460), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n479), .B1(new_n977), .B2(new_n508), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n973), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n476), .A2(G40), .A3(new_n484), .A4(new_n485), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT110), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n981), .A2(new_n982), .A3(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n723), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT109), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n783), .B(new_n789), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n723), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n984), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT111), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n824), .A2(new_n828), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n783), .A2(G2067), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n824), .A2(new_n828), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n998), .B2(new_n994), .ZN(new_n999));
  NOR2_X1   g574(.A1(G290), .A2(G1986), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n983), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT48), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n993), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n985), .B(KEYINPUT46), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n988), .A2(new_n723), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n991), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n997), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  AND4_X1   g584(.A1(G40), .A2(new_n476), .A3(new_n484), .A4(new_n485), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n981), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1971), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT112), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT50), .B1(new_n511), .B2(new_n973), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT50), .B(new_n973), .C1(new_n976), .C2(new_n978), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1010), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1015), .B(new_n1017), .C1(G2090), .C2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(G166), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(G8), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n982), .A2(new_n979), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n1026), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT114), .B1(new_n797), .B2(G1976), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n797), .A2(KEYINPUT114), .A3(G1976), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  NAND2_X1  g612(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n528), .A2(new_n580), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1039), .B2(new_n579), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(KEYINPUT116), .B2(KEYINPUT49), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT115), .B(G1981), .Z(new_n1042));
  AOI211_X1 g617(.A(new_n579), .B(new_n1042), .C1(new_n581), .C2(new_n583), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1038), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1042), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n584), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n1040), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1047), .A3(new_n1032), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1037), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1029), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n979), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n982), .B1(new_n1056), .B2(new_n1019), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT119), .ZN(new_n1058));
  AOI21_X1  g633(.A(G2090), .B1(new_n1057), .B2(KEYINPUT119), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1058), .A2(new_n1059), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1054), .B1(new_n1060), .B2(new_n1026), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1030), .A2(new_n1053), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2084), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1011), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n511), .B2(new_n973), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n1066), .B2(new_n982), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n486), .A2(new_n981), .A3(new_n1068), .A4(G40), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1064), .B1(new_n1070), .B2(G1966), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(G8), .A3(G168), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1009), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT121), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1052), .A2(KEYINPUT117), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1037), .A2(new_n1048), .A3(new_n1076), .A4(new_n1051), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1022), .A2(G8), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1072), .B1(new_n1080), .B2(new_n1054), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(KEYINPUT63), .A3(new_n1030), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(new_n1009), .C1(new_n1062), .C2(new_n1072), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1074), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1048), .A2(new_n1049), .A3(new_n797), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1032), .B1(new_n1086), .B2(new_n1043), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1078), .B2(new_n1030), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT118), .B(new_n1087), .C1(new_n1078), .C2(new_n1030), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G299), .B(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1010), .A2(new_n981), .A3(new_n1011), .A4(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1098), .C1(G1956), .C2(new_n1057), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1021), .A2(new_n713), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1094), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1010), .A2(new_n989), .A3(new_n981), .A4(new_n1011), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n982), .B2(new_n979), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n554), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1098), .B1(G1956), .B2(new_n1057), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT122), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1098), .B(new_n1112), .C1(G1956), .C2(new_n1057), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1096), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1099), .A2(KEYINPUT61), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1103), .B(new_n1109), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT123), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1096), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1113), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1112), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1103), .A4(new_n1109), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1021), .A2(new_n842), .B1(new_n789), .B2(new_n1031), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n598), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n598), .B1(new_n1126), .B2(KEYINPUT60), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1127), .A2(new_n1128), .B1(KEYINPUT60), .B2(new_n1126), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1117), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1100), .A2(new_n598), .A3(new_n1126), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1114), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(G2078), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1070), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1021), .A2(new_n705), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1134), .B1(new_n1012), .B2(G2078), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1136), .A2(KEYINPUT125), .A3(new_n1137), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G301), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1010), .A2(new_n1135), .A3(new_n981), .A4(new_n1011), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1141), .A2(G171), .A3(new_n1145), .A4(new_n1137), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(KEYINPUT54), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(G171), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1141), .A2(G301), .A3(new_n1145), .A4(new_n1137), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(KEYINPUT126), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(KEYINPUT126), .B2(new_n1150), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n1155));
  OAI211_X1 g730(.A(G168), .B(new_n1064), .C1(new_n1070), .C2(G1966), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G8), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1071), .A2(G286), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT51), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1156), .B2(G8), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1155), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1071), .B2(G286), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1157), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1167), .A2(KEYINPUT124), .A3(new_n1163), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1133), .A2(new_n1154), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1148), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1161), .A2(new_n1155), .A3(new_n1164), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT124), .B1(new_n1167), .B2(new_n1163), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1175), .A3(KEYINPUT62), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1062), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1093), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(G290), .A2(G1986), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n983), .B1(new_n1181), .B2(new_n1000), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n993), .A2(new_n1182), .A3(new_n999), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1008), .B1(new_n1180), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g759(.A1(new_n650), .A2(G319), .A3(new_n663), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1187));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1188));
  NAND4_X1  g762(.A1(new_n650), .A2(new_n1188), .A3(G319), .A4(new_n663), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1190), .A2(new_n915), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n959), .A3(new_n872), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1192), .A2(KEYINPUT43), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n958), .A2(new_n968), .A3(new_n964), .ZN(new_n1194));
  AOI211_X1 g768(.A(G229), .B(new_n1191), .C1(new_n1193), .C2(new_n1194), .ZN(G308));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  NAND4_X1  g770(.A1(new_n1196), .A2(new_n685), .A3(new_n915), .A4(new_n1190), .ZN(G225));
endmodule


