//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n468), .A2(G136), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT67), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n469), .B1(new_n466), .B2(new_n467), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(G162));
  NAND3_X1  g057(.A1(new_n461), .A2(G138), .A3(new_n469), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n476), .A2(G126), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n489), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n489), .B2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(G2104), .B(new_n488), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G88), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(G50), .A3(G543), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT70), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT70), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(G303));
  INV_X1    g084(.A(G303), .ZN(G166));
  NAND2_X1  g085(.A1(new_n500), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n496), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT72), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT73), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n499), .A2(KEYINPUT71), .A3(G63), .A4(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n514), .A2(new_n515), .B1(new_n497), .B2(new_n498), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT74), .B(G89), .Z(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n519), .A2(new_n522), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT76), .B(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(G651), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n536), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n518), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n526), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT77), .B(G81), .Z(new_n548));
  AOI22_X1  g123(.A1(new_n547), .A2(G651), .B1(new_n530), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n507), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n526), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n561), .A2(KEYINPUT78), .A3(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n500), .A2(G53), .A3(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n516), .A2(new_n566), .A3(G53), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n567), .B1(G91), .B2(new_n530), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  NAND3_X1  g144(.A1(new_n499), .A2(new_n500), .A3(G87), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n497), .A2(new_n571), .A3(new_n498), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n500), .A2(G49), .A3(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT79), .ZN(G288));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n497), .B2(new_n498), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT80), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(G73), .A3(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n499), .A2(new_n500), .A3(G86), .ZN(new_n585));
  AND2_X1   g160(.A1(KEYINPUT6), .A2(G651), .ZN(new_n586));
  NOR2_X1   g161(.A1(KEYINPUT6), .A2(G651), .ZN(new_n587));
  OAI211_X1 g162(.A(G48), .B(G543), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n518), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n526), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT81), .B(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n593), .A2(G651), .B1(new_n530), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n499), .A2(new_n500), .A3(G92), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n518), .A2(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n507), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G868), .ZN(G284));
  XOR2_X1   g180(.A(G284), .B(KEYINPUT82), .Z(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n476), .A2(G123), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT83), .Z(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G135), .B2(new_n468), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n461), .A2(new_n470), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(G2096), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n625), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G1341), .ZN(new_n642));
  INV_X1    g217(.A(G1348), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G1341), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G1348), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n651), .B1(new_n644), .B2(new_n647), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2084), .B(G2090), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  OR2_X1    g236(.A1(new_n656), .A2(KEYINPUT85), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(KEYINPUT85), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n658), .C2(new_n659), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(KEYINPUT86), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(KEYINPUT86), .ZN(new_n666));
  INV_X1    g241(.A(new_n658), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n659), .B(KEYINPUT17), .Z(new_n668));
  OAI211_X1 g243(.A(new_n665), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n657), .A3(new_n667), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT87), .B(G2096), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n683), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n687), .C1(new_n681), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n697));
  NOR2_X1   g272(.A1(G29), .A2(G35), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G162), .B2(G29), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT29), .B(G2090), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G4), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n604), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(new_n643), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(G20), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT23), .Z(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G299), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1956), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n701), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n468), .A2(G139), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n461), .A2(G127), .ZN(new_n715));
  NAND2_X1  g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n469), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(G33), .ZN(new_n721));
  INV_X1    g296(.A(G2072), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n702), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n702), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1966), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(new_n722), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT99), .B(G28), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(new_n719), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n623), .B2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n702), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n550), .B2(new_n702), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1341), .ZN(new_n738));
  OR4_X1    g313(.A1(new_n723), .A2(new_n726), .A3(new_n735), .A4(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n470), .A2(G105), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n740), .B(new_n742), .C1(G141), .C2(new_n468), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n476), .A2(G129), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT98), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(new_n719), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n719), .B2(G32), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n719), .B1(new_n752), .B2(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G160), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2084), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n749), .A2(new_n750), .ZN(new_n758));
  NOR2_X1   g333(.A1(G5), .A2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G301), .B2(new_n702), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n751), .A2(new_n757), .A3(new_n758), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n468), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n476), .A2(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n469), .A2(G116), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n719), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2067), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n719), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n719), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(G2078), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n761), .A2(new_n762), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n777), .B(new_n778), .C1(G2078), .C2(new_n776), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n710), .A2(new_n739), .A3(new_n764), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n702), .A2(G24), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G290), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT89), .B(G1986), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n468), .A2(G131), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n476), .A2(G119), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n469), .A2(G107), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G25), .B(new_n790), .S(G29), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT35), .B(G1991), .Z(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n785), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G6), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G16), .ZN(new_n797));
  AOI211_X1 g372(.A(KEYINPUT90), .B(new_n797), .C1(G305), .C2(G16), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n580), .A2(new_n582), .ZN(new_n800));
  OAI21_X1  g375(.A(G61), .B1(new_n524), .B2(new_n525), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n507), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n525), .A2(new_n524), .B1(new_n586), .B2(new_n587), .ZN(new_n803));
  INV_X1    g378(.A(G86), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n588), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(G16), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n797), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n799), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT32), .B(G1981), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT91), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n798), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n530), .A2(G86), .B1(new_n516), .B2(G48), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n702), .B1(new_n813), .B2(new_n584), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT90), .B1(new_n814), .B2(new_n797), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n806), .A2(new_n799), .A3(new_n807), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n508), .B(G16), .C1(new_n503), .C2(new_n504), .ZN(new_n819));
  OR2_X1    g394(.A1(G16), .A2(G22), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT92), .B(G1971), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n821), .B1(new_n819), .B2(new_n820), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT93), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n819), .A2(new_n820), .ZN(new_n825));
  INV_X1    g400(.A(new_n821), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT93), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n575), .A2(G16), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n702), .A2(G23), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n833), .ZN(new_n835));
  AOI211_X1 g410(.A(KEYINPUT33), .B(new_n835), .C1(new_n575), .C2(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(G1976), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n516), .A2(G49), .B1(new_n572), .B2(G651), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n702), .B1(new_n838), .B2(new_n570), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT33), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  INV_X1    g415(.A(G1976), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n832), .A2(new_n831), .A3(new_n833), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n818), .A2(new_n824), .A3(new_n830), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n795), .B1(new_n845), .B2(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT94), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n795), .B(new_n848), .C1(new_n845), .C2(KEYINPUT34), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n845), .A2(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT95), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n845), .A2(new_n854), .A3(KEYINPUT34), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND4_X1   g431(.A1(KEYINPUT97), .A2(new_n850), .A3(new_n851), .A4(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n847), .A2(new_n849), .B1(new_n853), .B2(new_n855), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT97), .B1(new_n858), .B2(new_n851), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT96), .B1(new_n858), .B2(new_n851), .ZN(new_n861));
  INV_X1    g436(.A(new_n849), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n815), .A2(new_n816), .A3(new_n810), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n811), .B1(new_n798), .B2(new_n808), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n844), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT34), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n824), .A4(new_n830), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n848), .B1(new_n867), .B2(new_n795), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n854), .B1(new_n845), .B2(KEYINPUT34), .ZN(new_n869));
  INV_X1    g444(.A(new_n855), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n862), .A2(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT36), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n861), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n697), .B(new_n781), .C1(new_n860), .C2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n871), .B2(KEYINPUT36), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n858), .A2(KEYINPUT97), .A3(new_n851), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n858), .A2(KEYINPUT96), .A3(new_n851), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n871), .B2(KEYINPUT36), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT101), .B1(new_n881), .B2(new_n780), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n875), .A2(new_n882), .ZN(G311));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n780), .ZN(G150));
  AOI22_X1  g459(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n885));
  INV_X1    g460(.A(G93), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n885), .A2(new_n507), .B1(new_n886), .B2(new_n803), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(G55), .B2(new_n518), .ZN(new_n888));
  INV_X1    g463(.A(G860), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT37), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n603), .A2(new_n611), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n550), .A2(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n544), .A2(new_n549), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n518), .A2(G55), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n897), .B2(new_n887), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n894), .B(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n889), .B1(new_n900), .B2(KEYINPUT39), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT103), .Z(G145));
  XNOR2_X1  g479(.A(G162), .B(G160), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n623), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n714), .A2(KEYINPUT104), .A3(new_n717), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n746), .B(new_n907), .Z(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(new_n769), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n769), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n493), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n476), .A2(G130), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n469), .A2(G118), .ZN(new_n914));
  OAI21_X1  g489(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(G142), .B2(new_n468), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n627), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n790), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n909), .A2(G164), .A3(new_n910), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n912), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(KEYINPUT105), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n912), .A2(new_n924), .A3(new_n919), .A4(new_n920), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n906), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n906), .A2(new_n921), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n922), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(G395));
  OAI21_X1  g507(.A(new_n607), .B1(new_n897), .B2(new_n887), .ZN(new_n933));
  XNOR2_X1  g508(.A(G303), .B(G290), .ZN(new_n934));
  XNOR2_X1  g509(.A(G305), .B(new_n575), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n603), .A2(G299), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n603), .A2(G299), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT41), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n944), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n942), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n942), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n899), .B(new_n613), .ZN(new_n952));
  MUX2_X1   g527(.A(new_n949), .B(new_n951), .S(new_n952), .Z(new_n953));
  NAND2_X1  g528(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT106), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n941), .A2(KEYINPUT108), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n939), .A3(new_n940), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n953), .A2(KEYINPUT108), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n933), .B1(new_n961), .B2(new_n607), .ZN(G295));
  OAI21_X1  g537(.A(new_n933), .B1(new_n961), .B2(new_n607), .ZN(G331));
  AND3_X1   g538(.A1(new_n895), .A2(G286), .A3(new_n898), .ZN(new_n964));
  AOI21_X1  g539(.A(G286), .B1(new_n895), .B2(new_n898), .ZN(new_n965));
  OAI21_X1  g540(.A(G301), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n899), .A2(G168), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n895), .A2(G286), .A3(new_n898), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(G171), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n951), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n949), .A2(new_n966), .A3(new_n969), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n936), .A4(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n974), .A2(new_n927), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n936), .A3(new_n973), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n949), .A2(KEYINPUT110), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n966), .B(new_n969), .C1(new_n979), .C2(new_n945), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n971), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n936), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n975), .A2(new_n977), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n971), .A2(new_n973), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n982), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n977), .A2(new_n987), .A3(new_n927), .A4(new_n974), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n985), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n975), .A2(new_n992), .A3(new_n977), .A4(new_n983), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g571(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n991), .C2(new_n993), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(G397));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n493), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n465), .A2(G40), .A3(new_n471), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n493), .A2(KEYINPUT112), .A3(new_n999), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(G1996), .A3(new_n746), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1009));
  INV_X1    g584(.A(G2067), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n769), .B(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n746), .B2(G1996), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1008), .A2(new_n1009), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n790), .A2(new_n793), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n793), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1006), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G290), .B(G1986), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1006), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n493), .B2(new_n999), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1004), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(G2078), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n493), .A2(new_n1028), .A3(new_n999), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1004), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n762), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1032), .A2(new_n1022), .A3(new_n1003), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1021), .A2(G2078), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1026), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1020), .B1(new_n1036), .B2(G171), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1024), .A2(new_n1034), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT122), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1005), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1044), .B2(new_n1003), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2078), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1033), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1048), .A2(new_n1021), .B1(new_n1030), .B2(new_n762), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(G301), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1037), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1046), .A2(new_n1020), .A3(new_n1049), .A4(G301), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT124), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1037), .A2(new_n1050), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1053), .A4(new_n1052), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(G166), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1022), .A2(new_n1003), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1971), .B1(new_n1066), .B2(new_n1024), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT114), .B(G2090), .Z(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1030), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n493), .A2(new_n1028), .A3(new_n999), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1028), .B1(new_n493), .B2(new_n999), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1003), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1067), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n1077));
  OAI21_X1  g652(.A(G8), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(KEYINPUT117), .B(new_n1067), .C1(new_n1071), .C2(new_n1075), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1065), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1049), .A2(G301), .A3(new_n1035), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1045), .B2(new_n1040), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT54), .B(new_n1081), .C1(new_n1083), .C2(G301), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G305), .A2(G1981), .ZN(new_n1086));
  INV_X1    g661(.A(G1981), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n813), .A2(new_n1087), .A3(new_n584), .ZN(new_n1088));
  OR2_X1    g663(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(new_n1061), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n838), .A2(G1976), .A3(new_n570), .ZN(new_n1095));
  OAI211_X1 g670(.A(G8), .B(new_n1095), .C1(new_n1000), .C2(new_n1003), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1092), .A2(new_n1094), .B1(KEYINPUT52), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n841), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1085), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1085), .A3(new_n1099), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1030), .A2(new_n1069), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1067), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1061), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1101), .A2(new_n1102), .B1(new_n1105), .B2(new_n1064), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1027), .A2(new_n1004), .A3(new_n756), .A4(new_n1029), .ZN(new_n1107));
  OAI211_X1 g682(.A(G168), .B(new_n1107), .C1(new_n1033), .C2(G1966), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  INV_X1    g684(.A(G1966), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1025), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G168), .B1(new_n1111), .B2(new_n1107), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT51), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1108), .A2(new_n1114), .A3(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AND4_X1   g691(.A1(new_n1080), .A2(new_n1084), .A3(new_n1106), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1059), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1023), .A2(new_n1004), .A3(new_n1024), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n563), .A2(new_n1121), .A3(new_n568), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n563), .B2(new_n568), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1120), .B(new_n1125), .C1(new_n1074), .C2(G1956), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1120), .B1(new_n1074), .B2(G1956), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1956), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1030), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(KEYINPUT119), .A3(new_n1125), .A4(new_n1120), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1125), .B1(new_n1133), .B2(new_n1120), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1140), .A2(new_n1128), .A3(KEYINPUT120), .A4(new_n1134), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT61), .B1(new_n1131), .B2(new_n1126), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT58), .B(G1341), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1025), .A2(G1996), .B1(new_n1093), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n550), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT121), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1142), .A2(new_n1152), .A3(new_n1149), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1030), .A2(new_n643), .B1(new_n1010), .B2(new_n1093), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT60), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(new_n604), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(KEYINPUT60), .B2(new_n1154), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1151), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1154), .A2(new_n603), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1126), .B1(new_n1159), .B2(new_n1138), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1118), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1092), .A2(G1976), .A3(G288), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1088), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1094), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1064), .B(G8), .C1(new_n1067), .C2(new_n1103), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1061), .B(G286), .C1(new_n1111), .C2(new_n1107), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1080), .A2(new_n1106), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1065), .B1(new_n1104), .B2(new_n1061), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1165), .A4(new_n1168), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1167), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1113), .A2(new_n1177), .A3(new_n1115), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1036), .A2(G171), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1097), .A2(new_n1085), .A3(new_n1099), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1165), .B1(new_n1182), .B2(new_n1100), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1068), .B1(new_n1074), .B2(KEYINPUT116), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1030), .A2(new_n1070), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1184), .A2(new_n1185), .B1(G1971), .B2(new_n1033), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT117), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(G8), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1183), .B1(new_n1189), .B2(new_n1065), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1176), .B1(new_n1181), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1180), .B1(new_n1116), .B2(KEYINPUT62), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1113), .A2(new_n1177), .A3(new_n1115), .ZN(new_n1193));
  AND4_X1   g768(.A1(new_n1176), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1175), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1019), .B1(new_n1161), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1006), .ZN(new_n1197));
  OR3_X1    g772(.A1(new_n1197), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT46), .B1(new_n1197), .B2(G1996), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n747), .A2(new_n1011), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n1199), .B1(new_n1006), .B2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT47), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1017), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT126), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1197), .A2(G1986), .A3(G290), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1206), .B(KEYINPUT48), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(G2067), .B2(new_n769), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1202), .B(new_n1208), .C1(new_n1006), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1196), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g787(.A(new_n459), .B1(new_n675), .B2(new_n676), .ZN(new_n1214));
  OAI211_X1 g788(.A(KEYINPUT127), .B(new_n1214), .C1(new_n653), .C2(new_n654), .ZN(new_n1215));
  AND2_X1   g789(.A1(new_n1215), .A2(new_n695), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1214), .B1(new_n653), .B2(new_n654), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g793(.A(new_n1216), .B(new_n1219), .C1(new_n926), .C2(new_n929), .ZN(new_n1220));
  INV_X1    g794(.A(new_n994), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n1220), .A2(new_n1221), .ZN(G308));
  OR2_X1    g796(.A1(new_n1220), .A2(new_n1221), .ZN(G225));
endmodule


