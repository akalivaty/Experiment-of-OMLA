//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n215));
  XNOR2_X1  g0015(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n209), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT1), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n227));
  AND3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n210), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n216), .B(new_n221), .C1(new_n222), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(new_n222), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n243), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT81), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G257), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT80), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n263), .A2(KEYINPUT80), .A3(G257), .A4(new_n253), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n254), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G303), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(G264), .A3(G1698), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n258), .A2(new_n264), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n219), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT66), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G1), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT5), .B(G41), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n277), .A2(G274), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT5), .A2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT5), .A2(G41), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n277), .A2(new_n285), .A3(G270), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n273), .A2(G179), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G116), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n219), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n208), .A2(G33), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G116), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G283), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n209), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G97), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n306), .B2(new_n260), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n293), .A2(new_n219), .B1(G20), .B2(new_n298), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n300), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT77), .B(G97), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT20), .B(new_n308), .C1(new_n312), .C2(new_n302), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n299), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n252), .B1(new_n289), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(new_n299), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n287), .B1(new_n268), .B2(new_n272), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT81), .A4(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n273), .A2(new_n288), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(new_n318), .A3(G169), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT21), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n322), .A2(new_n318), .A3(KEYINPUT21), .A4(G169), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n233), .A2(G1698), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G226), .B2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n330), .B2(new_n265), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n272), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(G41), .ZN(new_n334));
  AOI21_X1  g0134(.A(G1), .B1(new_n334), .B2(new_n278), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n277), .A2(G274), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n335), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n277), .A2(new_n337), .A3(G238), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n332), .A2(new_n333), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n219), .B1(new_n274), .B2(new_n270), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n335), .B1(new_n342), .B2(new_n276), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n331), .A2(new_n272), .B1(new_n343), .B2(G238), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(KEYINPUT72), .A3(new_n333), .A4(new_n336), .ZN(new_n345));
  NOR2_X1   g0145(.A1(G226), .A2(G1698), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n233), .B2(G1698), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n263), .B1(G33), .B2(G97), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n336), .B(new_n338), .C1(new_n348), .C2(new_n271), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n341), .A2(new_n345), .A3(G190), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n339), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G200), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT73), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n290), .B2(G68), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n246), .A2(G20), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n209), .A2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n209), .A2(new_n260), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n357), .B1(new_n358), .B2(new_n202), .C1(new_n244), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT11), .B1(new_n360), .B2(new_n294), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n208), .A2(G20), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n295), .A2(G68), .A3(new_n290), .A4(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n351), .A2(new_n353), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n343), .A2(G226), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n336), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(G1698), .B1(new_n261), .B2(new_n262), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G222), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n265), .A2(G77), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G1698), .B1(new_n254), .B2(new_n255), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT67), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT67), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n263), .A2(new_n378), .A3(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n375), .B1(G223), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n371), .B1(new_n381), .B2(new_n271), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G200), .ZN(new_n383));
  OAI211_X1 g0183(.A(G190), .B(new_n371), .C1(new_n381), .C2(new_n271), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n244), .B1(new_n208), .B2(G20), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n386), .A2(new_n219), .A3(new_n293), .A4(new_n290), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n208), .A2(new_n244), .A3(G13), .A4(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT68), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(KEYINPUT68), .A3(new_n388), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n209), .A2(new_n260), .A3(G150), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT8), .B(G58), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n392), .B1(new_n201), .B2(new_n209), .C1(new_n393), .C2(new_n358), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n390), .A2(new_n391), .B1(new_n294), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT9), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n294), .ZN(new_n398));
  INV_X1    g0198(.A(new_n391), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n389), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT9), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n400), .B2(new_n402), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT10), .B1(new_n397), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n384), .A2(new_n385), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT70), .B1(new_n395), .B2(KEYINPUT9), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n403), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n382), .A2(G200), .B1(KEYINPUT9), .B2(new_n395), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT10), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n408), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n290), .A2(new_n219), .A3(new_n293), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n364), .A2(G77), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n415), .A2(new_n416), .B1(G77), .B2(new_n290), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G20), .A2(G77), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n418), .B1(new_n419), .B2(new_n358), .C1(new_n359), .C2(new_n393), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n420), .B2(new_n294), .ZN(new_n421));
  OAI211_X1 g0221(.A(G232), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT69), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n422), .A2(new_n423), .B1(new_n265), .B2(G107), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n372), .A2(KEYINPUT69), .A3(G232), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G238), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n377), .B2(new_n379), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n272), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n343), .A2(G244), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n336), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n421), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n380), .A2(G238), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n425), .A3(new_n424), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n437), .B2(new_n272), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n429), .A2(new_n432), .A3(G190), .ZN(new_n442));
  INV_X1    g0242(.A(G200), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n421), .B(new_n442), .C1(new_n438), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n380), .A2(G223), .ZN(new_n445));
  INV_X1    g0245(.A(new_n375), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n271), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n370), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n439), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n400), .C1(G169), .C2(new_n448), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n414), .A2(new_n441), .A3(new_n444), .A4(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n439), .B1(new_n349), .B2(KEYINPUT13), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n341), .A2(new_n452), .A3(new_n345), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT74), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n341), .A2(new_n452), .A3(new_n345), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT14), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n352), .B2(G169), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT14), .B(new_n434), .C1(new_n350), .C2(new_n339), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n366), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n277), .A2(new_n337), .A3(G232), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G87), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT76), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(KEYINPUT76), .A2(G33), .A3(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G223), .A2(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G226), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G1698), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n263), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n336), .B(new_n464), .C1(new_n473), .C2(new_n271), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n434), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(G179), .B2(new_n474), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n261), .A2(new_n209), .A3(new_n262), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT7), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n262), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n246), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G58), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n246), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G58), .A2(G68), .ZN(new_n484));
  OAI21_X1  g0284(.A(G20), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G159), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n359), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT75), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT16), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT75), .B(new_n490), .C1(new_n481), .C2(new_n487), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n294), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n393), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n364), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n494), .A2(new_n415), .B1(new_n290), .B2(new_n493), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n476), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT18), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n295), .B1(new_n488), .B2(KEYINPUT16), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n495), .B1(new_n500), .B2(new_n491), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT18), .B1(new_n501), .B2(new_n476), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n474), .A2(new_n443), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n471), .A2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G223), .B2(G1698), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n467), .B(new_n468), .C1(new_n506), .C2(new_n265), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n272), .ZN(new_n508));
  INV_X1    g0308(.A(G190), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n336), .A4(new_n464), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n492), .A2(new_n496), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT17), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n501), .A2(KEYINPUT17), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n503), .A2(new_n516), .ZN(new_n517));
  AND4_X1   g0317(.A1(new_n368), .A2(new_n451), .A3(new_n463), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n322), .A2(G200), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n314), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n314), .B(new_n519), .C1(new_n319), .C2(new_n443), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n319), .A2(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT83), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n319), .A2(new_n443), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT82), .B1(new_n526), .B2(new_n318), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n523), .A4(new_n522), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n372), .A2(KEYINPUT4), .A3(G244), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n301), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n272), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n277), .A2(new_n285), .A3(G257), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n281), .A2(new_n538), .A3(KEYINPUT78), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT78), .B1(new_n281), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n290), .A2(G97), .ZN(new_n543));
  INV_X1    g0343(.A(new_n297), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n479), .A2(new_n480), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G107), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n303), .B2(new_n305), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT6), .B1(new_n206), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G20), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n548), .B(new_n553), .C1(new_n202), .C2(new_n359), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n546), .B1(new_n554), .B2(new_n294), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n281), .A2(new_n538), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n536), .B2(new_n272), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G190), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n542), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n419), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n290), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n209), .B1(new_n328), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n205), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n306), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n311), .B2(new_n358), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n263), .A2(new_n209), .A3(G68), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n561), .B1(new_n569), .B2(new_n294), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n544), .A2(new_n560), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  INV_X1    g0373(.A(G244), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n573), .C1(new_n376), .C2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G250), .B1(new_n208), .B2(G45), .ZN(new_n576));
  INV_X1    g0376(.A(G274), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n279), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n575), .A2(new_n272), .B1(new_n277), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n570), .A2(new_n571), .B1(new_n579), .B2(new_n439), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G169), .B2(new_n579), .ZN(new_n581));
  INV_X1    g0381(.A(new_n556), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n537), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n434), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n553), .B1(new_n202), .B2(new_n359), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n205), .B1(new_n479), .B2(new_n480), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n294), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n545), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n537), .B(new_n439), .C1(new_n540), .C2(new_n539), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n297), .A2(new_n564), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n561), .B(new_n591), .C1(new_n569), .C2(new_n294), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n579), .A2(KEYINPUT79), .A3(G190), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT79), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n575), .A2(new_n272), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n578), .A2(new_n277), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n597), .B2(G200), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n595), .A2(G190), .A3(new_n596), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n593), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n559), .A2(new_n581), .A3(new_n590), .A4(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n209), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n263), .A2(new_n604), .A3(new_n209), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n573), .A2(G20), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT23), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n209), .B2(G107), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT24), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n606), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n294), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n277), .A2(new_n285), .A3(G264), .ZN(new_n618));
  OAI211_X1 g0418(.A(G250), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n619));
  OAI211_X1 g0419(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G33), .A2(G294), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT84), .A4(new_n621), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n272), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n281), .B(new_n618), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G200), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT25), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n290), .B2(G107), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n290), .A2(new_n629), .A3(G107), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n544), .A2(G107), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n622), .A2(new_n623), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n272), .A3(new_n625), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(G190), .A3(new_n281), .A4(new_n618), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n617), .A2(new_n628), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n627), .A2(new_n434), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n439), .A3(new_n281), .A4(new_n618), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n295), .B1(new_n613), .B2(new_n615), .ZN(new_n640));
  INV_X1    g0440(.A(new_n633), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n601), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n327), .A2(new_n518), .A3(new_n530), .A4(new_n644), .ZN(G372));
  INV_X1    g0445(.A(KEYINPUT85), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n575), .A2(new_n646), .A3(new_n272), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n575), .B2(new_n272), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n596), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n434), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n580), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n434), .A2(new_n583), .B1(new_n587), .B2(new_n545), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n600), .A2(new_n581), .A3(new_n653), .A4(new_n589), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n654), .B2(KEYINPUT26), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n591), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n570), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n599), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n649), .A2(G200), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n656), .A2(new_n657), .A3(new_n651), .A4(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n321), .A2(new_n642), .A3(new_n325), .A4(new_n326), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n661), .A2(new_n660), .B1(new_n650), .B2(new_n580), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n637), .A3(new_n590), .A4(new_n559), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n655), .B(new_n663), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n518), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n450), .ZN(new_n669));
  INV_X1    g0469(.A(new_n463), .ZN(new_n670));
  INV_X1    g0470(.A(new_n368), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n441), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n502), .B(new_n499), .C1(new_n673), .C2(new_n516), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT86), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n414), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n407), .A2(KEYINPUT86), .A3(new_n413), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n669), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n668), .A2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT27), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n208), .A3(new_n209), .A4(G13), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(G213), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n640), .B2(new_n641), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n637), .A2(new_n642), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT89), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  INV_X1    g0493(.A(new_n642), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n688), .ZN(new_n695));
  INV_X1    g0495(.A(new_n688), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n530), .B(new_n327), .C1(new_n314), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n327), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n318), .A3(new_n688), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT88), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT88), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n703), .A3(G330), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n695), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n327), .A2(new_n688), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n692), .A2(new_n706), .A3(new_n693), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n694), .A2(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n705), .A2(new_n709), .ZN(G399));
  NOR3_X1   g0510(.A1(new_n306), .A2(G116), .A3(new_n565), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT90), .Z(new_n712));
  NOR2_X1   g0512(.A1(new_n212), .A2(G41), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n712), .A2(new_n208), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n218), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT91), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT28), .Z(new_n717));
  NOR2_X1   g0517(.A1(new_n664), .A2(new_n666), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n651), .A3(new_n663), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n696), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n667), .A2(KEYINPUT93), .A3(new_n696), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n651), .B1(new_n654), .B2(KEYINPUT26), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n657), .B1(new_n665), .B2(new_n656), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n642), .A2(new_n321), .A3(new_n325), .A4(new_n326), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n559), .A2(new_n590), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n637), .A4(new_n665), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n688), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n644), .A2(new_n530), .A3(new_n327), .A4(new_n696), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n541), .A2(new_n627), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n541), .A2(new_n627), .A3(KEYINPUT92), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n649), .A2(new_n439), .A3(new_n322), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n557), .A2(new_n618), .A3(new_n635), .A4(new_n579), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(new_n289), .ZN(new_n745));
  INV_X1    g0545(.A(new_n289), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n537), .A2(new_n579), .A3(new_n582), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n635), .A2(new_n618), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT30), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n688), .B1(new_n742), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(KEYINPUT31), .B(new_n688), .C1(new_n742), .C2(new_n750), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n736), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n735), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n717), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n219), .B1(G20), .B2(new_n434), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n212), .A2(new_n263), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n278), .B2(new_n218), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n250), .B2(new_n278), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n212), .A2(new_n265), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G355), .B1(new_n298), .B2(new_n212), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n765), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n209), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n439), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n263), .B1(new_n775), .B2(new_n202), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n209), .A2(new_n439), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n509), .A3(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n246), .B1(new_n779), .B2(new_n244), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n209), .A2(new_n509), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n774), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n776), .B(new_n780), .C1(G58), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n443), .A2(G179), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n781), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n773), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n784), .B1(new_n564), .B2(new_n787), .C1(new_n205), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n439), .A2(new_n443), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n773), .ZN(new_n793));
  OR3_X1    g0593(.A1(new_n793), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT32), .B1(new_n793), .B2(new_n486), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n209), .B1(new_n792), .B2(G190), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n795), .C1(new_n204), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n793), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n788), .C1(new_n801), .C2(new_n787), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n775), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n263), .B(new_n804), .C1(G322), .C2(new_n783), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  INV_X1    g0606(.A(new_n778), .ZN(new_n807));
  INV_X1    g0607(.A(new_n779), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(G326), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n805), .B(new_n809), .C1(new_n810), .C2(new_n796), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n789), .A2(new_n797), .B1(new_n802), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n772), .B1(new_n812), .B2(new_n763), .ZN(new_n813));
  INV_X1    g0613(.A(new_n762), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n700), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n702), .B(new_n704), .C1(G330), .C2(new_n700), .ZN(new_n816));
  INV_X1    g0616(.A(new_n713), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n211), .A2(G20), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n208), .B1(new_n818), .B2(G45), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n817), .A2(KEYINPUT94), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT94), .ZN(new_n821));
  INV_X1    g0621(.A(new_n819), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n713), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  MUX2_X1   g0624(.A(new_n815), .B(new_n816), .S(new_n824), .Z(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT97), .ZN(G396));
  OR3_X1    g0626(.A1(new_n421), .A2(new_n686), .A3(new_n687), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n444), .A2(new_n827), .B1(new_n440), .B2(new_n435), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n435), .A2(new_n440), .A3(new_n696), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT100), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n442), .A2(new_n421), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n443), .B1(new_n429), .B2(new_n432), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n441), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n435), .A2(new_n440), .A3(new_n696), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n667), .A2(new_n838), .A3(new_n696), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n723), .A2(new_n725), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(new_n756), .ZN(new_n842));
  INV_X1    g0642(.A(new_n824), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n841), .B2(new_n756), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n763), .A2(new_n760), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n843), .B1(G77), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n788), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G68), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n793), .ZN(new_n852));
  INV_X1    g0652(.A(new_n787), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n265), .B(new_n852), .C1(G50), .C2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n482), .B2(new_n796), .ZN(new_n855));
  INV_X1    g0655(.A(new_n775), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n783), .B1(new_n856), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n779), .C1(new_n859), .C2(new_n778), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  OAI22_X1  g0661(.A1(new_n796), .A2(new_n204), .B1(new_n810), .B2(new_n782), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT99), .Z(new_n863));
  OAI21_X1  g0663(.A(new_n265), .B1(new_n787), .B2(new_n205), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT98), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n798), .A2(G311), .B1(new_n849), .B2(G87), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(KEYINPUT98), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n779), .A2(new_n801), .B1(new_n775), .B2(new_n298), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G283), .B2(new_n807), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n855), .A2(new_n861), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n848), .B1(new_n871), .B2(new_n763), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n761), .B2(new_n838), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT101), .Z(new_n874));
  NOR2_X1   g0674(.A1(new_n845), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  OR2_X1    g0676(.A1(new_n550), .A2(new_n552), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n220), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OAI211_X1 g0681(.A(new_n218), .B(G77), .C1(new_n482), .C2(new_n246), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n208), .B(G13), .C1(new_n882), .C2(new_n245), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n492), .A2(new_n496), .ZN(new_n885));
  INV_X1    g0685(.A(new_n476), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n686), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .A4(new_n512), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  AOI221_X4 g0692(.A(new_n495), .B1(new_n504), .B2(new_n510), .C1(new_n500), .C2(new_n491), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n497), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n890), .A4(new_n889), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n512), .B1(new_n501), .B2(new_n476), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n501), .A2(new_n686), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n892), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n503), .B2(new_n516), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n891), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n901), .A3(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n366), .A2(new_n688), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n463), .A2(new_n368), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n366), .B(new_n688), .C1(new_n462), .C2(new_n671), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n909), .A2(new_n910), .B1(new_n837), .B2(new_n830), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n911), .A2(new_n755), .A3(KEYINPUT40), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n905), .A2(new_n901), .A3(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n905), .B2(new_n901), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n755), .B(new_n911), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n907), .A2(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n518), .A3(new_n755), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n518), .B2(new_n755), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n900), .B2(new_n901), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n905), .A2(new_n901), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n903), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n924), .A2(new_n670), .A3(new_n696), .A4(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n909), .A2(new_n910), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n839), .B2(new_n836), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n906), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n930), .A2(new_n931), .B1(new_n503), .B2(new_n686), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n726), .A2(new_n518), .A3(new_n734), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n679), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n921), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n208), .B2(new_n818), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n921), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n884), .B1(new_n938), .B2(new_n939), .ZN(G367));
  NOR2_X1   g0740(.A1(new_n590), .A2(new_n696), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT104), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n731), .B1(new_n555), .B2(new_n696), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n705), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT103), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n696), .A2(new_n592), .ZN(new_n947));
  MUX2_X1   g0747(.A(new_n665), .B(new_n652), .S(new_n947), .Z(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n944), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(new_n707), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n590), .B1(new_n954), .B2(new_n642), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n955), .A2(KEYINPUT42), .B1(new_n956), .B2(new_n696), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n957), .A2(new_n958), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n953), .B(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n713), .B(KEYINPUT41), .Z(new_n961));
  AOI21_X1  g0761(.A(new_n944), .B1(new_n708), .B2(new_n707), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(KEYINPUT44), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n707), .A2(new_n944), .A3(new_n708), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n963), .A2(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT105), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n705), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT106), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n969), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT106), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(new_n977), .A3(new_n971), .A4(new_n705), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n702), .A2(new_n704), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n695), .B1(new_n327), .B2(new_n688), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n707), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n758), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n975), .A2(new_n705), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n974), .A2(new_n978), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n961), .B1(new_n986), .B2(new_n758), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT107), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n819), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(KEYINPUT107), .B(new_n961), .C1(new_n986), .C2(new_n758), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n960), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n239), .A2(new_n766), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n764), .B1(new_n213), .B2(new_n419), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n263), .B1(new_n775), .B2(new_n244), .C1(new_n778), .C2(new_n486), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n793), .A2(new_n858), .B1(new_n787), .B2(new_n482), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G77), .C2(new_n849), .ZN(new_n996));
  INV_X1    g0796(.A(G143), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n779), .A2(new_n997), .B1(new_n782), .B2(new_n859), .ZN(new_n998));
  INV_X1    g0798(.A(new_n796), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(G68), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n265), .B1(new_n788), .B2(new_n311), .C1(new_n793), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT108), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G303), .A2(new_n783), .B1(new_n856), .B2(G283), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n810), .B2(new_n778), .C1(new_n803), .C2(new_n779), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n999), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n853), .A2(G116), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT46), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1003), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  INV_X1    g0816(.A(new_n763), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n843), .B1(new_n992), .B2(new_n993), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n814), .C2(new_n948), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n991), .A2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n982), .A2(new_n822), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n695), .A2(new_n762), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n796), .A2(new_n800), .B1(new_n810), .B2(new_n787), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n782), .A2(new_n1004), .B1(new_n775), .B2(new_n801), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT111), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(KEYINPUT111), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n807), .A2(G311), .B1(new_n808), .B2(G322), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1025), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n263), .B1(new_n798), .B2(G326), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n298), .C2(new_n788), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT49), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n787), .A2(new_n202), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G97), .B2(new_n849), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n859), .B2(new_n793), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n796), .A2(new_n419), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n263), .B1(new_n775), .B2(new_n246), .C1(new_n244), .C2(new_n782), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n486), .A2(new_n779), .B1(new_n778), .B2(new_n393), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n763), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n236), .A2(new_n278), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1047), .A2(new_n766), .B1(new_n712), .B2(new_n770), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n393), .A2(G50), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT50), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n278), .B1(new_n246), .B2(new_n202), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1051), .B(new_n712), .C1(new_n1050), .C2(new_n1049), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1048), .A2(new_n1052), .B1(G107), .B2(new_n213), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n824), .B1(new_n1053), .B2(new_n764), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1024), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n983), .A2(new_n713), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n982), .A2(new_n758), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1023), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(G393));
  XOR2_X1   g0858(.A(new_n969), .B(new_n705), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n817), .B1(new_n1059), .B2(new_n983), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n986), .A2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1059), .A2(new_n819), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n764), .B1(new_n213), .B2(new_n311), .C1(new_n243), .C2(new_n767), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(new_n843), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n793), .A2(new_n997), .B1(new_n787), .B2(new_n246), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n265), .B(new_n1065), .C1(G87), .C2(new_n849), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n778), .A2(new_n244), .B1(new_n775), .B2(new_n393), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n808), .A2(G150), .B1(new_n783), .B2(G159), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1070), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n999), .A2(G77), .B1(new_n1074), .B2(new_n1071), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1067), .A2(new_n1068), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT52), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n779), .A2(new_n1004), .B1(new_n782), .B2(new_n803), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n999), .A2(G116), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n265), .B1(new_n775), .B2(new_n810), .C1(new_n778), .C2(new_n801), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n849), .B2(G107), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n798), .A2(G322), .B1(new_n853), .B2(G283), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1078), .A2(new_n1077), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1064), .B1(new_n944), .B2(new_n814), .C1(new_n1086), .C2(new_n1017), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1061), .A2(new_n1062), .A3(new_n1087), .ZN(G390));
  OAI21_X1  g0888(.A(new_n265), .B1(new_n787), .B2(new_n564), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT118), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n778), .A2(new_n205), .B1(new_n775), .B2(new_n311), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n999), .A2(G77), .B1(KEYINPUT117), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(KEYINPUT117), .B2(new_n1091), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n808), .A2(G283), .B1(new_n783), .B2(G116), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n850), .B(new_n1094), .C1(new_n810), .C2(new_n793), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n798), .A2(G125), .B1(new_n849), .B2(G50), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n775), .A2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n265), .B(new_n1099), .C1(G132), .C2(new_n783), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n807), .A2(G137), .B1(new_n808), .B2(G128), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G159), .B2(new_n999), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n787), .A2(new_n859), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1090), .A2(new_n1096), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n843), .B1(new_n493), .B2(new_n847), .C1(new_n1106), .C2(new_n1017), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n924), .A2(new_n927), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n760), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n839), .A2(new_n836), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n909), .A2(new_n910), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n670), .A2(new_n696), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n924), .A2(new_n927), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n755), .A2(G330), .A3(new_n838), .A4(new_n1112), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(KEYINPUT115), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n733), .A2(new_n838), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n929), .B1(new_n1119), .B2(new_n836), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n923), .B2(new_n913), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1115), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1108), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1117), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1110), .B1(new_n1128), .B2(new_n819), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n757), .A2(new_n518), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n934), .A2(new_n679), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n755), .A2(G330), .A3(new_n838), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n929), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1116), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1111), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n829), .B1(new_n733), .B2(new_n838), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1116), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1132), .A2(KEYINPUT116), .A3(new_n929), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1131), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1127), .B2(new_n1123), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n817), .B1(new_n1128), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1129), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n395), .A2(new_n686), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n678), .B2(new_n450), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n407), .A2(KEYINPUT86), .A3(new_n413), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT86), .B1(new_n407), .B2(new_n413), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n450), .B(new_n1151), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n450), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1150), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1155), .A3(new_n1148), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n760), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n843), .B1(G50), .B2(new_n847), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n788), .A2(new_n482), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1039), .B(new_n1165), .C1(G283), .C2(new_n798), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n334), .B(new_n265), .C1(new_n775), .C2(new_n419), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n778), .A2(new_n204), .B1(new_n779), .B2(new_n298), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(G107), .C2(new_n783), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1166), .B(new_n1169), .C1(new_n246), .C2(new_n796), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n265), .A2(new_n334), .ZN(new_n1172));
  AOI21_X1  g0972(.A(G50), .B1(new_n260), .B2(new_n334), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1170), .A2(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n778), .A2(new_n851), .ZN(new_n1175));
  INV_X1    g0975(.A(G128), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n782), .A2(new_n1176), .B1(new_n775), .B2(new_n858), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G125), .C2(new_n808), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n859), .B2(new_n796), .C1(new_n787), .C2(new_n1098), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n260), .B(new_n334), .C1(new_n788), .C2(new_n486), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G124), .B2(new_n798), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1174), .B1(new_n1171), .B2(new_n1170), .C1(new_n1180), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1164), .B1(new_n1185), .B2(new_n763), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1163), .A2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT119), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n907), .A2(new_n912), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n915), .A2(new_n916), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(G330), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n1162), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1161), .B1(new_n917), .B2(G330), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n933), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1162), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n928), .A2(new_n932), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n917), .A2(G330), .A3(new_n1161), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n819), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1188), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1196), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1118), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1125), .A2(new_n1126), .A3(new_n1117), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1141), .A2(new_n1135), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1131), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(KEYINPUT120), .B(new_n713), .C1(new_n1203), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1208), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1210), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1131), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1143), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT120), .B1(new_n1217), .B2(new_n713), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1200), .B1(new_n1213), .B2(new_n1218), .ZN(G375));
  INV_X1    g1019(.A(new_n1207), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1131), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n961), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1144), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n929), .A2(new_n760), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT121), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n847), .A2(G68), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G77), .A2(new_n849), .B1(new_n853), .B2(G97), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n801), .B2(new_n793), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n265), .B1(new_n775), .B2(new_n205), .C1(new_n800), .C2(new_n782), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n778), .A2(new_n298), .B1(new_n779), .B2(new_n810), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1228), .A2(new_n1042), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT122), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1165), .B1(G159), .B2(new_n853), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n999), .A2(G50), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n263), .B1(new_n782), .B2(new_n858), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n851), .A2(new_n779), .B1(new_n778), .B2(new_n1098), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(G150), .C2(new_n856), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n798), .A2(G128), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1234), .A2(new_n1235), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1232), .A2(KEYINPUT122), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1233), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n824), .B(new_n1226), .C1(new_n1242), .C2(new_n763), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1207), .A2(new_n822), .B1(new_n1225), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1223), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT123), .ZN(G381));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n875), .A3(new_n1146), .A4(new_n1248), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(G387), .A2(G375), .A3(G381), .A4(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT124), .Z(G407));
  INV_X1    g1051(.A(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(G375), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G378), .A2(G343), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G407), .A2(new_n1255), .ZN(G409));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  NAND3_X1  g1057(.A1(new_n991), .A2(new_n1021), .A3(new_n1247), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1247), .B1(new_n991), .B2(new_n1021), .ZN(new_n1260));
  OAI211_X1 g1060(.A(KEYINPUT126), .B(new_n1257), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(G390), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1258), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1252), .A2(G343), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G378), .B(new_n1200), .C1(new_n1213), .C2(new_n1218), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1216), .B(new_n1222), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1270), .B(new_n1187), .C1(new_n1211), .C2(new_n819), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1187), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT125), .B1(new_n1199), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1146), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1267), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1221), .B1(new_n1277), .B2(new_n1142), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1220), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n713), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1244), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n875), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(G384), .A3(new_n1244), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1276), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1268), .A2(new_n1275), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1267), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT127), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1289), .B(new_n1267), .C1(new_n1268), .C2(new_n1275), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1267), .A2(G2897), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1282), .A2(new_n1283), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1266), .B1(new_n1293), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1297), .B2(new_n1276), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT63), .B1(new_n1276), .B2(new_n1284), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1303), .A2(new_n1306), .A3(new_n1261), .A4(new_n1265), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1302), .A2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1146), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1268), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1284), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1266), .B(new_n1311), .ZN(G402));
endmodule


