//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G71gat), .ZN(new_n202));
  INV_X1    g001(.A(G78gat), .ZN(new_n203));
  OAI211_X1 g002(.A(new_n202), .B(new_n203), .C1(KEYINPUT97), .C2(KEYINPUT9), .ZN(new_n204));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n207), .B2(KEYINPUT97), .ZN(new_n208));
  OR2_X1    g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT96), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT96), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(KEYINPUT9), .A3(new_n210), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT95), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT95), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G71gat), .B2(G78gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n217), .A3(new_n219), .A4(new_n205), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(G1gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT93), .ZN(new_n230));
  AOI21_X1  g029(.A(G8gat), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n231), .B(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n222), .B2(new_n221), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT98), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n227), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G155gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G183gat), .B(G211gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n238), .B(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(G232gat), .A2(G233gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT41), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT99), .ZN(new_n246));
  XNOR2_X1  g045(.A(G134gat), .B(G162gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT88), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n254), .A2(KEYINPUT89), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n254), .A2(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258));
  OR2_X1    g057(.A1(G43gat), .A2(G50gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(G43gat), .A2(G50gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OR3_X1    g060(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT92), .B(G50gat), .Z(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G43gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT91), .B(G43gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G50gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n258), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT90), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n261), .A2(new_n269), .B1(G29gat), .B2(G36gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n262), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n268), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n263), .A2(KEYINPUT17), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(G99gat), .A2(G106gat), .ZN(new_n278));
  INV_X1    g077(.A(G85gat), .ZN(new_n279));
  INV_X1    g078(.A(G92gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(KEYINPUT8), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G99gat), .B(G106gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT7), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n279), .B2(new_n280), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n281), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT100), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(new_n282), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n287), .A3(new_n286), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n288), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n288), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n274), .A2(new_n294), .B1(KEYINPUT41), .B2(new_n244), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G190gat), .B(G218gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n296), .A2(new_n297), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n249), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n296), .A2(new_n297), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n248), .A3(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n243), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n291), .A2(new_n286), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n307), .A2(KEYINPUT101), .A3(new_n220), .A4(new_n215), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT101), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n286), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n221), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n221), .A3(new_n288), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n308), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n215), .A2(new_n220), .A3(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT102), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n294), .A2(KEYINPUT102), .A3(new_n315), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G230gat), .A2(G233gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n308), .A2(new_n312), .A3(new_n311), .ZN(new_n323));
  INV_X1    g122(.A(new_n321), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G120gat), .B(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  NAND3_X1  g128(.A1(new_n322), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT103), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n325), .B1(new_n321), .B2(new_n320), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT103), .A3(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n333), .A2(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n306), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT65), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(G169gat), .A3(G176gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT66), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT25), .B1(new_n345), .B2(KEYINPUT23), .ZN(new_n349));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT24), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n349), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n344), .A2(new_n358), .A3(new_n346), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361));
  INV_X1    g160(.A(G183gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(KEYINPUT24), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n363), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n350), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT64), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G169gat), .ZN(new_n370));
  INV_X1    g169(.A(G176gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n344), .A2(new_n346), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n361), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(KEYINPUT28), .A3(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n345), .B(KEYINPUT26), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n384), .A2(new_n344), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n360), .A2(new_n376), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G134gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G127gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n226), .A2(G134gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT1), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT67), .ZN(new_n392));
  INV_X1    g191(.A(G120gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(G113gat), .ZN(new_n394));
  INV_X1    g193(.A(G113gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n394), .B(new_n396), .C1(new_n395), .C2(G120gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n395), .A2(G120gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n393), .A2(G113gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n391), .A2(new_n397), .B1(new_n401), .B2(new_n390), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT69), .B1(new_n386), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n385), .ZN(new_n404));
  INV_X1    g203(.A(new_n349), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n364), .B2(new_n355), .ZN(new_n406));
  AOI221_X4 g205(.A(KEYINPUT66), .B1(new_n345), .B2(KEYINPUT23), .C1(new_n341), .C2(new_n343), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n358), .B1(new_n344), .B2(new_n346), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n344), .A2(new_n346), .A3(new_n374), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n354), .A2(new_n367), .A3(new_n366), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT25), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n404), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT69), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n397), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n401), .A2(new_n390), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n360), .A2(new_n376), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n402), .A3(new_n404), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT68), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n386), .A2(new_n423), .A3(new_n402), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT34), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n403), .A2(new_n418), .B1(new_n422), .B2(new_n424), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n427), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT33), .B1(new_n426), .B2(new_n428), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT70), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(new_n202), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(G99gat), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n429), .B(new_n432), .C1(new_n433), .C2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n430), .B2(new_n427), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n431), .B1(new_n430), .B2(new_n427), .ZN(new_n442));
  AND4_X1   g241(.A1(new_n431), .A2(new_n419), .A3(new_n425), .A4(new_n427), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n441), .B(new_n437), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n428), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT32), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n439), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n439), .B2(new_n444), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G78gat), .B(G106gat), .Z(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT82), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(G50gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  INV_X1    g257(.A(G148gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G141gat), .ZN(new_n460));
  INV_X1    g259(.A(G141gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G148gat), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT76), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G155gat), .B(G162gat), .ZN(new_n464));
  INV_X1    g263(.A(G155gat), .ZN(new_n465));
  INV_X1    g264(.A(G162gat), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT2), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n463), .B2(new_n467), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G211gat), .B(G218gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT72), .ZN(new_n473));
  INV_X1    g272(.A(G197gat), .ZN(new_n474));
  INV_X1    g273(.A(G204gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G197gat), .A2(G204gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT22), .ZN(new_n478));
  NAND2_X1  g277(.A1(G211gat), .A2(G218gat), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n481), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n471), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n460), .A2(new_n462), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT76), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n467), .ZN(new_n490));
  INV_X1    g289(.A(new_n464), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n486), .A3(new_n468), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n482), .A2(new_n483), .B1(new_n493), .B2(new_n484), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT83), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G22gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT83), .B(G22gat), .C1(new_n487), .C2(new_n494), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n497), .B2(new_n500), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n457), .B(new_n458), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n501), .A2(new_n502), .A3(new_n457), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n450), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT3), .B1(new_n469), .B2(new_n470), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n493), .A3(new_n417), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n492), .A2(new_n415), .A3(new_n468), .A4(new_n416), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n471), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n516));
  NAND4_X1  g315(.A1(new_n514), .A2(KEYINPUT79), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT79), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n509), .A2(new_n513), .A3(new_n512), .A4(new_n515), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n492), .A2(new_n468), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n417), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n510), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n417), .A3(KEYINPUT77), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(G225gat), .A3(G233gat), .A4(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n517), .A2(new_n521), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G1gat), .B(G29gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT0), .ZN(new_n531));
  XNOR2_X1  g330(.A(G57gat), .B(G85gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  AOI21_X1  g332(.A(KEYINPUT6), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT80), .B1(new_n529), .B2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n521), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n522), .A2(new_n528), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT80), .ZN(new_n539));
  INV_X1    g338(.A(new_n533), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n534), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(KEYINPUT6), .A3(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n482), .A2(new_n483), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g345(.A1(G226gat), .A2(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n420), .A2(KEYINPUT73), .A3(new_n404), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT73), .B1(new_n420), .B2(new_n404), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n546), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT73), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n413), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n386), .A2(KEYINPUT73), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n413), .A2(new_n484), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT74), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n545), .B(new_n551), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n554), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n548), .A2(KEYINPUT29), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n545), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n386), .A2(new_n548), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G8gat), .B(G36gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G64gat), .B(G92gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT75), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n568), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n558), .B2(new_n564), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT75), .B1(new_n574), .B2(KEYINPUT30), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n565), .A2(KEYINPUT30), .A3(new_n568), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n564), .A3(new_n573), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n544), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT35), .B1(new_n507), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n575), .B2(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n538), .A2(new_n540), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n534), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT35), .B1(new_n585), .B2(new_n543), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n450), .A2(new_n506), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n505), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n503), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n559), .A2(new_n560), .B1(new_n548), .B2(new_n386), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT37), .B1(new_n592), .B2(new_n562), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n547), .B1(new_n386), .B2(KEYINPUT29), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n546), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n545), .B1(new_n597), .B2(new_n551), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n591), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n573), .A2(KEYINPUT37), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n578), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n536), .A2(new_n533), .A3(new_n537), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT6), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n529), .A2(new_n533), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n569), .B(new_n543), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n578), .A2(new_n600), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n565), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT38), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n590), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT87), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n514), .A2(KEYINPUT39), .A3(new_n515), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n526), .A2(new_n527), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n515), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n616), .B(KEYINPUT39), .C1(new_n515), .C2(new_n514), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n617), .A3(new_n533), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT86), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n621), .A3(new_n619), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n618), .B2(new_n619), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n584), .B(new_n620), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n613), .B1(new_n583), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n574), .A2(KEYINPUT75), .A3(KEYINPUT30), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n579), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n584), .B1(new_n619), .B2(new_n618), .ZN(new_n630));
  INV_X1    g429(.A(new_n624), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n631), .B2(new_n622), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(KEYINPUT87), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n439), .A2(new_n444), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n446), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n439), .A2(new_n444), .A3(new_n447), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n448), .B2(new_n449), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n640), .A2(new_n642), .B1(new_n580), .B2(new_n590), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT85), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n634), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n580), .A2(new_n590), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT85), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n588), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G197gat), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT11), .B(G169gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT13), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n235), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n274), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n235), .A2(new_n273), .A3(new_n263), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n276), .A2(new_n235), .A3(new_n277), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n656), .A3(new_n660), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT18), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n663), .A2(KEYINPUT18), .A3(new_n656), .A4(new_n660), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n655), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n655), .A3(new_n667), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n650), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT94), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n650), .A2(KEYINPUT94), .A3(new_n671), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n339), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n544), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  INV_X1    g479(.A(new_n671), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n648), .A2(KEYINPUT85), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n643), .A2(new_n644), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n634), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n673), .B(new_n681), .C1(new_n684), .C2(new_n588), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT94), .B1(new_n650), .B2(new_n671), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n629), .B(new_n338), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT16), .B(G8gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n680), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n691), .B(new_n680), .C1(new_n687), .C2(new_n688), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n687), .A2(new_n680), .A3(new_n688), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(G8gat), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n690), .A2(new_n692), .A3(new_n693), .A4(new_n694), .ZN(G1325gat));
  OAI21_X1  g494(.A(new_n338), .B1(new_n685), .B2(new_n686), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n646), .A2(KEYINPUT105), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n642), .A2(new_n640), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G15gat), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n450), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(G15gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n676), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(KEYINPUT106), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n676), .A2(new_n590), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n305), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n650), .A2(new_n715), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n634), .A2(new_n643), .B1(new_n581), .B2(new_n587), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(new_n305), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n243), .A2(new_n337), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n681), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n713), .B1(new_n723), .B2(new_n544), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n719), .A2(KEYINPUT107), .A3(new_n677), .A4(new_n722), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(G29gat), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n721), .A2(new_n305), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n674), .B2(new_n675), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n544), .A2(G29gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n730), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n726), .A2(new_n733), .A3(new_n734), .ZN(G1328gat));
  NOR2_X1   g534(.A1(new_n583), .A2(G36gat), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n727), .B(new_n736), .C1(new_n685), .C2(new_n686), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n723), .B2(new_n583), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(G1329gat));
  INV_X1    g542(.A(new_n700), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n716), .A2(new_n744), .A3(new_n718), .A4(new_n722), .ZN(new_n745));
  INV_X1    g544(.A(new_n266), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n745), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n702), .A2(new_n746), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n727), .B(new_n751), .C1(new_n685), .C2(new_n686), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n723), .B2(new_n646), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1330gat));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n716), .A2(new_n590), .A3(new_n718), .A4(new_n722), .ZN(new_n760));
  INV_X1    g559(.A(new_n264), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n506), .A2(new_n761), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n727), .B(new_n763), .C1(new_n685), .C2(new_n686), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(KEYINPUT110), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n729), .B2(new_n763), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n759), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n264), .B1(new_n760), .B2(KEYINPUT111), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT111), .B2(new_n760), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(KEYINPUT48), .A3(new_n764), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1331gat));
  INV_X1    g571(.A(new_n337), .ZN(new_n773));
  NOR4_X1   g572(.A1(new_n717), .A2(new_n671), .A3(new_n306), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n677), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g575(.A(new_n583), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT112), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n779), .B(new_n780), .Z(G1333gat));
  AOI21_X1  g580(.A(new_n202), .B1(new_n774), .B2(new_n744), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n702), .A2(G71gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n774), .A2(new_n590), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g586(.A1(new_n717), .A2(new_n305), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n243), .A2(new_n671), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n788), .A2(KEYINPUT51), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n279), .A3(new_n677), .A4(new_n337), .ZN(new_n793));
  INV_X1    g592(.A(new_n789), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n773), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n719), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n544), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1336gat));
  NOR3_X1   g597(.A1(new_n583), .A2(G92gat), .A3(new_n773), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT113), .Z(new_n800));
  NAND3_X1  g599(.A1(new_n719), .A2(new_n629), .A3(new_n795), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n792), .A2(new_n800), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n801), .A2(G92gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n799), .B1(new_n790), .B2(new_n791), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n803), .ZN(new_n806));
  OAI22_X1  g605(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n806), .ZN(G1337gat));
  NOR2_X1   g606(.A1(new_n702), .A2(G99gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n337), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT114), .B1(new_n796), .B2(new_n700), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G99gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n796), .A2(KEYINPUT114), .A3(new_n700), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(G1338gat));
  NOR2_X1   g612(.A1(new_n506), .A2(G106gat), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n337), .B(new_n814), .C1(new_n790), .C2(new_n791), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n716), .A2(new_n590), .A3(new_n718), .A4(new_n795), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n314), .A2(new_n318), .A3(new_n324), .A4(new_n319), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n322), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n329), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n320), .A2(new_n824), .A3(new_n321), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n664), .A2(new_n665), .ZN(new_n829));
  INV_X1    g628(.A(new_n662), .ZN(new_n830));
  AND4_X1   g629(.A1(new_n655), .A2(new_n829), .A3(new_n830), .A4(new_n667), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n831), .B2(new_n668), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n823), .A4(new_n825), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n335), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n335), .A2(KEYINPUT115), .A3(new_n833), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n656), .B1(new_n663), .B2(new_n660), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n660), .A2(new_n661), .A3(new_n658), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n654), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n337), .A2(new_n670), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n305), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n335), .A2(KEYINPUT115), .A3(new_n833), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT115), .B1(new_n335), .B2(new_n833), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n304), .A2(new_n670), .A3(new_n841), .A4(new_n828), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n243), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n306), .A2(new_n671), .A3(new_n337), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n820), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n243), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n671), .B(new_n828), .C1(new_n845), .C2(new_n846), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n304), .B1(new_n854), .B2(new_n842), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n847), .A2(new_n848), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n851), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT116), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n702), .A2(new_n544), .A3(new_n629), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n506), .A3(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n395), .A3(new_n681), .ZN(new_n863));
  INV_X1    g662(.A(new_n507), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n852), .A2(new_n859), .A3(new_n677), .A4(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n629), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n671), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n863), .B1(new_n395), .B2(new_n869), .ZN(G1340gat));
  NAND2_X1  g669(.A1(new_n337), .A2(new_n393), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT118), .Z(new_n872));
  NAND3_X1  g671(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G120gat), .B1(new_n862), .B2(new_n773), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1341gat));
  NAND4_X1  g676(.A1(new_n867), .A2(new_n868), .A3(new_n226), .A4(new_n243), .ZN(new_n878));
  OAI21_X1  g677(.A(G127gat), .B1(new_n862), .B2(new_n853), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  NAND4_X1  g679(.A1(new_n867), .A2(new_n868), .A3(new_n387), .A4(new_n304), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n862), .B2(new_n305), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1343gat));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n852), .A2(new_n859), .A3(new_n886), .A4(new_n590), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n629), .A2(new_n544), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n646), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n842), .B1(new_n832), .B2(new_n834), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n305), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n243), .B1(new_n849), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n590), .B1(new_n892), .B2(new_n851), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n671), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n860), .A2(new_n897), .A3(new_n677), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n852), .A2(new_n859), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT120), .B1(new_n899), .B2(new_n544), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n744), .A2(new_n629), .A3(new_n506), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n671), .A2(new_n461), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n896), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n895), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n895), .A2(new_n906), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n907), .A2(new_n908), .A3(new_n461), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n902), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n905), .B1(new_n909), .B2(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n646), .A2(new_n337), .A3(new_n888), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n852), .A2(new_n859), .A3(KEYINPUT57), .A4(new_n590), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n886), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n459), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n887), .A2(new_n894), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n773), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(KEYINPUT59), .A3(new_n459), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n337), .A2(new_n459), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n921), .A2(new_n924), .B1(new_n902), .B2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n922), .B2(new_n853), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n243), .A2(new_n465), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n902), .B2(new_n928), .ZN(G1346gat));
  NOR3_X1   g728(.A1(new_n922), .A2(new_n466), .A3(new_n305), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n902), .A2(new_n305), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n466), .ZN(G1347gat));
  NOR3_X1   g731(.A1(new_n702), .A2(new_n677), .A3(new_n583), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n860), .A2(new_n506), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n370), .A3(new_n681), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n507), .A2(new_n583), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT123), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n899), .A2(new_n677), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n671), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n935), .A2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n934), .B2(new_n773), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n371), .A3(new_n337), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n934), .B2(new_n853), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n243), .A2(new_n377), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n938), .A2(new_n945), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g746(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n934), .B2(new_n305), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT61), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n378), .A3(new_n304), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1351gat));
  AOI211_X1 g752(.A(new_n583), .B(new_n506), .C1(new_n697), .C2(new_n699), .ZN(new_n954));
  AND4_X1   g753(.A1(new_n544), .A2(new_n852), .A3(new_n859), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n671), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n700), .A2(new_n544), .A3(new_n629), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n915), .B2(new_n916), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n681), .A2(new_n474), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND4_X1  g759(.A1(new_n852), .A2(new_n859), .A3(new_n954), .A4(new_n544), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n773), .A2(G204gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT125), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n967));
  NOR4_X1   g766(.A1(new_n961), .A2(new_n967), .A3(KEYINPUT62), .A4(new_n963), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT62), .B1(new_n961), .B2(new_n963), .ZN(new_n970));
  AOI211_X1 g769(.A(new_n773), .B(new_n957), .C1(new_n915), .C2(new_n916), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n475), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT126), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n965), .A3(new_n962), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n967), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n964), .A2(KEYINPUT125), .A3(new_n965), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n958), .A2(new_n337), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G204gat), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n977), .A2(new_n978), .A3(new_n970), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n973), .A2(new_n981), .ZN(G1353gat));
  OR3_X1    g781(.A1(new_n961), .A2(G211gat), .A3(new_n853), .ZN(new_n983));
  OAI21_X1  g782(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n958), .B2(new_n243), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  INV_X1    g787(.A(G218gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n955), .A2(new_n989), .A3(new_n304), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n958), .A2(new_n304), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n990), .B1(new_n991), .B2(new_n989), .ZN(G1355gat));
endmodule


