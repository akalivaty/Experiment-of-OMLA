

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U324 ( .A(n344), .B(KEYINPUT32), .ZN(n345) );
  XNOR2_X1 U325 ( .A(n366), .B(KEYINPUT48), .ZN(n522) );
  INV_X1 U326 ( .A(n522), .ZN(n524) );
  XNOR2_X1 U327 ( .A(n346), .B(n345), .ZN(n349) );
  XOR2_X1 U328 ( .A(n354), .B(n353), .Z(n467) );
  XOR2_X1 U329 ( .A(KEYINPUT41), .B(n467), .Z(n543) );
  INV_X1 U330 ( .A(KEYINPUT123), .ZN(n448) );
  XOR2_X1 U331 ( .A(n553), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U332 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U333 ( .A(n451), .B(n450), .ZN(G1352GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n447) );
  XOR2_X1 U335 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n293) );
  XNOR2_X1 U336 ( .A(G92GAT), .B(KEYINPUT74), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n309) );
  XOR2_X1 U338 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n295) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n297) );
  XNOR2_X1 U341 ( .A(G36GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n296), .B(G218GAT), .ZN(n371) );
  XOR2_X1 U343 ( .A(n297), .B(n371), .Z(n303) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G43GAT), .Z(n299) );
  XNOR2_X1 U345 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n327) );
  XOR2_X1 U347 ( .A(KEYINPUT68), .B(G85GAT), .Z(n301) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n347) );
  XNOR2_X1 U350 ( .A(n327), .B(n347), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U352 ( .A(n304), .B(KEYINPUT10), .Z(n307) );
  XNOR2_X1 U353 ( .A(G50GAT), .B(KEYINPUT71), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n305), .B(G162GAT), .ZN(n425) );
  XNOR2_X1 U355 ( .A(G134GAT), .B(n425), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n568) );
  INV_X1 U358 ( .A(n568), .ZN(n463) );
  XOR2_X1 U359 ( .A(KEYINPUT75), .B(G211GAT), .Z(n311) );
  XNOR2_X1 U360 ( .A(G8GAT), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n369) );
  XOR2_X1 U362 ( .A(KEYINPUT76), .B(n369), .Z(n313) );
  NAND2_X1 U363 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U365 ( .A(n314), .B(G64GAT), .Z(n316) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G155GAT), .Z(n413) );
  XNOR2_X1 U367 ( .A(G127GAT), .B(n413), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U369 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n318) );
  XNOR2_X1 U370 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U372 ( .A(n320), .B(n319), .Z(n325) );
  XNOR2_X1 U373 ( .A(G15GAT), .B(G1GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n321), .B(KEYINPUT66), .ZN(n326) );
  XOR2_X1 U375 ( .A(KEYINPUT13), .B(G57GAT), .Z(n323) );
  XNOR2_X1 U376 ( .A(G71GAT), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n352) );
  XNOR2_X1 U378 ( .A(n326), .B(n352), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n577) );
  XNOR2_X1 U380 ( .A(n577), .B(KEYINPUT110), .ZN(n563) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n340) );
  XOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n329) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U385 ( .A(n330), .B(KEYINPUT30), .Z(n338) );
  XOR2_X1 U386 ( .A(G113GAT), .B(G36GAT), .Z(n332) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(G50GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U389 ( .A(G8GAT), .B(G141GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(G22GAT), .B(G197GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U394 ( .A(n340), .B(n339), .Z(n557) );
  INV_X1 U395 ( .A(n557), .ZN(n500) );
  XOR2_X1 U396 ( .A(KEYINPUT67), .B(G148GAT), .Z(n417) );
  XOR2_X1 U397 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n342) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n417), .B(n343), .Z(n346) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XOR2_X1 U402 ( .A(n347), .B(KEYINPUT69), .Z(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U404 ( .A(G64GAT), .B(G92GAT), .Z(n351) );
  XNOR2_X1 U405 ( .A(G176GAT), .B(G204GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n372) );
  XOR2_X1 U407 ( .A(n372), .B(n352), .Z(n353) );
  NOR2_X1 U408 ( .A1(n500), .A2(n543), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n355), .B(KEYINPUT46), .ZN(n356) );
  NOR2_X1 U410 ( .A1(n563), .A2(n356), .ZN(n357) );
  NAND2_X1 U411 ( .A1(n463), .A2(n357), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n358), .B(KEYINPUT47), .ZN(n365) );
  XOR2_X1 U413 ( .A(KEYINPUT36), .B(n463), .Z(n580) );
  NAND2_X1 U414 ( .A1(n580), .A2(n577), .ZN(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT111), .B(KEYINPUT45), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n359), .B(KEYINPUT64), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U418 ( .A1(n362), .A2(n467), .ZN(n363) );
  NOR2_X1 U419 ( .A1(n557), .A2(n363), .ZN(n364) );
  NOR2_X1 U420 ( .A1(n365), .A2(n364), .ZN(n366) );
  XOR2_X1 U421 ( .A(G197GAT), .B(KEYINPUT21), .Z(n412) );
  XOR2_X1 U422 ( .A(KEYINPUT94), .B(n412), .Z(n368) );
  NAND2_X1 U423 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U425 ( .A(n370), .B(n369), .Z(n374) );
  XNOR2_X1 U426 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U428 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n376) );
  XNOR2_X1 U429 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(n377), .ZN(n443) );
  INV_X1 U432 ( .A(n443), .ZN(n378) );
  XOR2_X1 U433 ( .A(n379), .B(n378), .Z(n472) );
  INV_X1 U434 ( .A(n472), .ZN(n516) );
  XNOR2_X1 U435 ( .A(KEYINPUT118), .B(n516), .ZN(n380) );
  NOR2_X1 U436 ( .A1(n522), .A2(n380), .ZN(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT54), .B(n381), .ZN(n405) );
  XOR2_X1 U438 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n383) );
  XNOR2_X1 U439 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n392) );
  XOR2_X1 U441 ( .A(KEYINPUT89), .B(KEYINPUT93), .Z(n390) );
  XOR2_X1 U442 ( .A(G127GAT), .B(G134GAT), .Z(n385) );
  XNOR2_X1 U443 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U445 ( .A(G113GAT), .B(n386), .Z(n431) );
  XOR2_X1 U446 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n388) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(KEYINPUT86), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n424) );
  XNOR2_X1 U449 ( .A(n431), .B(n424), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n404) );
  NAND2_X1 U452 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XOR2_X1 U453 ( .A(G57GAT), .B(G85GAT), .Z(n394) );
  XNOR2_X1 U454 ( .A(G148GAT), .B(G155GAT), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U456 ( .A(G29GAT), .B(G162GAT), .Z(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U459 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n400) );
  XNOR2_X1 U460 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U463 ( .A(n404), .B(n403), .Z(n469) );
  INV_X1 U464 ( .A(n469), .ZN(n513) );
  NAND2_X1 U465 ( .A1(n405), .A2(n513), .ZN(n552) );
  XOR2_X1 U466 ( .A(KEYINPUT24), .B(G78GAT), .Z(n407) );
  XNOR2_X1 U467 ( .A(G218GAT), .B(G106GAT), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT23), .B(G204GAT), .Z(n409) );
  XNOR2_X1 U470 ( .A(KEYINPUT88), .B(KEYINPUT85), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U472 ( .A(n411), .B(n410), .Z(n419) );
  XOR2_X1 U473 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U478 ( .A(G211GAT), .B(KEYINPUT22), .Z(n421) );
  XNOR2_X1 U479 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U481 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n553) );
  XOR2_X1 U484 ( .A(G71GAT), .B(KEYINPUT80), .Z(n429) );
  NAND2_X1 U485 ( .A1(G227GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n430), .B(G99GAT), .Z(n433) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT79), .B(KEYINPUT82), .Z(n435) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U493 ( .A(KEYINPUT20), .B(G176GAT), .Z(n437) );
  XNOR2_X1 U494 ( .A(G190GAT), .B(G183GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U496 ( .A(n439), .B(n438), .Z(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X2 U498 ( .A(n443), .B(n442), .Z(n556) );
  NAND2_X1 U499 ( .A1(n553), .A2(n556), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n444), .B(KEYINPUT26), .ZN(n539) );
  NOR2_X1 U501 ( .A1(n552), .A2(n539), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT122), .ZN(n581) );
  NAND2_X1 U503 ( .A1(n581), .A2(n557), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n451) );
  XNOR2_X1 U505 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n449) );
  INV_X1 U506 ( .A(n527), .ZN(n478) );
  XNOR2_X1 U507 ( .A(n516), .B(KEYINPUT27), .ZN(n456) );
  NOR2_X1 U508 ( .A1(n513), .A2(n456), .ZN(n523) );
  NAND2_X1 U509 ( .A1(n556), .A2(n523), .ZN(n452) );
  NOR2_X1 U510 ( .A1(n478), .A2(n452), .ZN(n462) );
  NOR2_X1 U511 ( .A1(n556), .A2(n516), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n553), .A2(n453), .ZN(n454) );
  XOR2_X1 U513 ( .A(n454), .B(KEYINPUT25), .Z(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT96), .B(n455), .Z(n459) );
  NOR2_X1 U515 ( .A1(n456), .A2(n539), .ZN(n457) );
  XNOR2_X1 U516 ( .A(KEYINPUT95), .B(n457), .ZN(n458) );
  AND2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U518 ( .A1(n460), .A2(n469), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n462), .A2(n461), .ZN(n483) );
  NAND2_X1 U520 ( .A1(n577), .A2(n463), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT78), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n465), .B(KEYINPUT16), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n483), .A2(n466), .ZN(n501) );
  INV_X1 U524 ( .A(n467), .ZN(n572) );
  NOR2_X1 U525 ( .A1(n500), .A2(n572), .ZN(n487) );
  NAND2_X1 U526 ( .A1(n501), .A2(n487), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT97), .ZN(n479) );
  NAND2_X1 U528 ( .A1(n469), .A2(n479), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n479), .A2(n472), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT98), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n477) );
  INV_X1 U535 ( .A(n556), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n479), .A2(n475), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  XOR2_X1 U538 ( .A(G22GAT), .B(KEYINPUT99), .Z(n481) );
  NAND2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1327GAT) );
  XNOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT101), .ZN(n490) );
  NOR2_X1 U543 ( .A1(n577), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT100), .B(n484), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n485), .A2(n580), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT37), .ZN(n512) );
  NAND2_X1 U547 ( .A1(n512), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT38), .B(n488), .ZN(n497) );
  NOR2_X1 U549 ( .A1(n513), .A2(n497), .ZN(n489) );
  XOR2_X1 U550 ( .A(n490), .B(n489), .Z(G1328GAT) );
  NOR2_X1 U551 ( .A1(n497), .A2(n516), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT102), .B(n491), .Z(n492) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n494) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n556), .A2(n497), .ZN(n495) );
  XOR2_X1 U558 ( .A(n496), .B(n495), .Z(G1330GAT) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n527), .A2(n497), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(n543), .B(KEYINPUT106), .Z(n559) );
  AND2_X1 U563 ( .A1(n500), .A2(n559), .ZN(n511) );
  NAND2_X1 U564 ( .A1(n511), .A2(n501), .ZN(n507) );
  NOR2_X1 U565 ( .A1(n513), .A2(n507), .ZN(n502) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n516), .A2(n507), .ZN(n504) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n556), .A2(n507), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  NOR2_X1 U573 ( .A1(n527), .A2(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n519) );
  NOR2_X1 U578 ( .A1(n513), .A2(n519), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n556), .A2(n519), .ZN(n518) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n527), .A2(n519), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(n520), .Z(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT112), .B(n525), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n556), .A2(n538), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(KEYINPUT113), .B(n528), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n557), .A2(n534), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U596 ( .A1(n534), .A2(n559), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U598 ( .A1(n563), .A2(n534), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n568), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT115), .B(n540), .ZN(n542) );
  INV_X1 U607 ( .A(n542), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n550), .A2(n557), .ZN(n541) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(n546), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n577), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n568), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT55), .ZN(n555) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n557), .A2(n569), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n569), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n569), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT119), .B(n567), .Z(n571) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n581), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n581), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

