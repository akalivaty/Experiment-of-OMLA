//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(G20), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n209), .A2(new_n220), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G150), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n248), .A2(G20), .A3(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n204), .B1(new_n221), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  AOI211_X1 g0055(.A(new_n249), .B(new_n251), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n226), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n204), .A3(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n203), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n262), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(G50), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT68), .B(G223), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(new_n278), .B1(G77), .B2(new_n275), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n281), .B(new_n282), .C1(new_n273), .C2(new_n274), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G222), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n272), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n272), .A3(G274), .ZN(new_n290));
  INV_X1    g0090(.A(G226), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n272), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G190), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n260), .A2(new_n269), .A3(new_n267), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n270), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(G200), .B1(new_n286), .B2(new_n294), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT71), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n298), .A2(new_n305), .A3(new_n301), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n295), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n268), .C1(G169), .C2(new_n295), .ZN(new_n310));
  INV_X1    g0110(.A(G244), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n290), .B1(new_n311), .B2(new_n293), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n284), .A2(G232), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n277), .A2(G238), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n275), .A2(G107), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n272), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n308), .B2(new_n318), .ZN(new_n320));
  INV_X1    g0120(.A(G77), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n203), .B2(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n263), .A2(new_n322), .B1(new_n321), .B2(new_n262), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT69), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n255), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G20), .A2(G33), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n253), .A2(new_n328), .B1(G20), .B2(G77), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n259), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI211_X1 g0132(.A(KEYINPUT70), .B(new_n259), .C1(new_n327), .C2(new_n329), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n320), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n318), .A2(G190), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n318), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n307), .A2(new_n310), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n328), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n342));
  INV_X1    g0142(.A(new_n255), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n321), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT11), .B1(new_n344), .B2(new_n258), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT75), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n347), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n345), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n266), .A2(KEYINPUT12), .A3(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT12), .B1(new_n266), .B2(G68), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n211), .B1(new_n203), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n352), .A2(new_n353), .B1(new_n263), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(G232), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(new_n283), .C2(new_n291), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n317), .ZN(new_n360));
  INV_X1    g0160(.A(new_n293), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n272), .A2(G274), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(G238), .A2(new_n361), .B1(new_n363), .B2(new_n289), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n360), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n360), .B2(new_n364), .ZN(new_n368));
  OAI21_X1  g0168(.A(G200), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n360), .A2(new_n364), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT13), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n366), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(G200), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n356), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n360), .A2(new_n364), .A3(KEYINPUT73), .A4(new_n365), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n372), .A3(G190), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n368), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n378), .A4(new_n379), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT14), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n373), .A2(new_n390), .A3(G169), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n378), .A2(new_n372), .A3(G179), .A4(new_n379), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n356), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n263), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n253), .A2(new_n264), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n397), .B1(new_n266), .B2(new_n253), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(G159), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n400), .A2(G20), .A3(G33), .ZN(new_n401));
  XNOR2_X1  g0201(.A(G58), .B(G68), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n399), .B(new_n401), .C1(G20), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT76), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n254), .ZN(new_n406));
  NAND2_X1  g0206(.A1(KEYINPUT3), .A2(G33), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n204), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n406), .A2(new_n410), .A3(new_n204), .A4(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n404), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G68), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n403), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n258), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT77), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(G68), .A3(new_n411), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n402), .A2(G20), .B1(G159), .B2(new_n328), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n421), .B2(new_n399), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT16), .B1(new_n419), .B2(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n418), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n398), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n272), .A2(G232), .A3(new_n292), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n290), .A2(new_n427), .A3(KEYINPUT78), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT78), .B1(new_n290), .B2(new_n427), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(G226), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  INV_X1    g0232(.A(G223), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n432), .C1(new_n283), .C2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(G179), .B1(new_n434), .B2(new_n317), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT79), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n290), .A2(new_n427), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n434), .B2(new_n317), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(G169), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n430), .A2(new_n435), .A3(KEYINPUT79), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT18), .B1(new_n426), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  INV_X1    g0246(.A(new_n398), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n416), .B(new_n258), .C1(new_n424), .C2(new_n418), .ZN(new_n448));
  INV_X1    g0248(.A(new_n425), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n430), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n434), .A2(new_n317), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT80), .A2(G190), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT80), .A2(G190), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n452), .A2(new_n457), .B1(G200), .B2(new_n440), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n423), .A2(new_n425), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(KEYINPUT17), .A3(new_n447), .A4(new_n458), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n444), .A2(new_n451), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n341), .A2(new_n395), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n326), .A2(new_n266), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n266), .B(new_n259), .C1(G1), .C2(new_n254), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n326), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n204), .B1(new_n471), .B2(new_n358), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT86), .ZN(new_n473));
  NOR3_X1   g0273(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT86), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n204), .C1(new_n471), .C2(new_n358), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n275), .A2(G20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n255), .A2(G97), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n479), .A2(G68), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n467), .B(new_n470), .C1(new_n482), .C2(new_n259), .ZN(new_n483));
  OAI211_X1 g0283(.A(G244), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G116), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n485), .C1(new_n283), .C2(new_n212), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n317), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n203), .A2(G45), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n272), .A2(G250), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n362), .B2(new_n488), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n486), .B2(new_n317), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n308), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G169), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n493), .B(new_n490), .C1(new_n317), .C2(new_n486), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT84), .B1(new_n487), .B2(new_n491), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n483), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n259), .B1(new_n478), .B2(new_n481), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n468), .A2(new_n213), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n503), .A2(new_n466), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(G190), .A3(new_n496), .ZN(new_n506));
  OAI21_X1  g0306(.A(G200), .B1(new_n499), .B2(new_n500), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n204), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT22), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n406), .A2(new_n407), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT22), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n204), .A4(G87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  OR3_X1    g0316(.A1(new_n485), .A2(KEYINPUT87), .A3(G20), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n204), .B2(G107), .ZN(new_n519));
  INV_X1    g0319(.A(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(KEYINPUT23), .A3(G20), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT87), .B1(new_n485), .B2(G20), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n516), .B1(new_n515), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n258), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n266), .B2(G107), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n266), .A2(new_n529), .A3(G107), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(new_n520), .B2(new_n468), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT5), .B(G41), .ZN(new_n535));
  INV_X1    g0335(.A(new_n488), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n537), .A2(G264), .A3(new_n272), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n512), .A2(G257), .A3(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G294), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(new_n540), .C1(new_n214), .C2(new_n283), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n317), .ZN(new_n542));
  INV_X1    g0342(.A(new_n537), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n363), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n542), .A2(new_n383), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(G200), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n528), .B(new_n534), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n541), .A2(new_n317), .ZN(new_n548));
  INV_X1    g0348(.A(new_n538), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n498), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n542), .A2(new_n308), .A3(new_n544), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n515), .A2(new_n524), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT24), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n259), .B1(new_n554), .B2(new_n525), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n551), .B(new_n552), .C1(new_n555), .C2(new_n533), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n547), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n263), .B(G116), .C1(G1), .C2(new_n254), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n262), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G283), .ZN(new_n561));
  INV_X1    g0361(.A(G97), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n204), .C1(G33), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(G20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n258), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n558), .B(new_n560), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n512), .A2(G264), .A3(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n275), .A2(G303), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n512), .A2(G257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n281), .A2(new_n282), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n317), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n317), .B1(new_n536), .B2(new_n535), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G270), .B1(new_n543), .B2(new_n363), .ZN(new_n578));
  INV_X1    g0378(.A(new_n456), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n576), .A2(new_n578), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n570), .B(new_n580), .C1(new_n581), .C2(new_n337), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n576), .A2(new_n578), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(G169), .A3(new_n569), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(G179), .A3(new_n569), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n569), .A3(KEYINPUT21), .A4(G169), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n582), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n509), .A2(new_n557), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n281), .A2(new_n282), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(KEYINPUT4), .A3(G244), .A4(new_n512), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n284), .A2(new_n594), .A3(KEYINPUT4), .A4(G244), .ZN(new_n595));
  INV_X1    g0395(.A(new_n561), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n277), .B2(G250), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n283), .B2(new_n311), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n593), .A2(new_n595), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n317), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n577), .A2(G257), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n544), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(KEYINPUT82), .A3(G200), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n328), .A2(G77), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT6), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n608), .A2(new_n562), .A3(G107), .ZN(new_n609));
  XNOR2_X1  g0409(.A(G97), .B(G107), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n607), .B1(new_n611), .B2(new_n204), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n409), .A2(G107), .A3(new_n411), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n258), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n266), .A2(G97), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n469), .B2(G97), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n603), .B1(new_n600), .B2(new_n317), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(G190), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT82), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n618), .B2(new_n337), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n606), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n308), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(new_n617), .C1(G169), .C2(new_n618), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n622), .A2(KEYINPUT83), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT83), .B1(new_n622), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n590), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n465), .A2(new_n627), .ZN(G372));
  NOR3_X1   g0428(.A1(new_n341), .A2(new_n395), .A3(new_n464), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n483), .B(new_n497), .C1(G169), .C2(new_n495), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n505), .B(new_n506), .C1(new_n337), .C2(new_n495), .ZN(new_n631));
  INV_X1    g0431(.A(new_n556), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n547), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n622), .A2(new_n624), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n509), .A2(new_n624), .A3(KEYINPUT88), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(new_n631), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n640), .B2(new_n624), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n502), .A2(new_n508), .ZN(new_n642));
  INV_X1    g0442(.A(new_n624), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n644), .A3(KEYINPUT88), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n461), .A2(new_n463), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n387), .A2(new_n335), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n394), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n444), .A2(new_n451), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n307), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n647), .A2(new_n310), .A3(new_n652), .ZN(G369));
  NAND3_X1  g0453(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n570), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n633), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n589), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n555), .A2(new_n533), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n660), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n557), .A2(new_n667), .B1(new_n556), .B2(new_n660), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n633), .A2(new_n660), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n557), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n632), .B2(new_n660), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(G399));
  NAND2_X1  g0473(.A1(new_n474), .A2(new_n559), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT89), .Z(new_n675));
  INV_X1    g0475(.A(new_n207), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n675), .A2(new_n677), .A3(new_n203), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n225), .B2(new_n677), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT28), .Z(new_n680));
  AOI21_X1  g0480(.A(new_n659), .B1(new_n639), .B2(new_n645), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n581), .A2(G179), .A3(new_n495), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n605), .A3(new_n550), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n576), .A2(new_n578), .A3(G179), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n548), .A2(new_n549), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n499), .A2(new_n500), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n618), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n691), .A2(KEYINPUT90), .A3(KEYINPUT30), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT30), .B1(new_n691), .B2(KEYINPUT90), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n684), .B(new_n686), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n627), .A2(KEYINPUT31), .B1(new_n659), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  INV_X1    g0496(.A(new_n686), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(KEYINPUT90), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n691), .A2(KEYINPUT90), .A3(KEYINPUT30), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n659), .A2(KEYINPUT31), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n696), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n686), .B1(new_n692), .B2(new_n693), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT91), .A3(KEYINPUT31), .A4(new_n659), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(G330), .B1(new_n695), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT26), .B1(new_n640), .B2(new_n624), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n642), .A2(new_n637), .A3(new_n643), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n660), .B1(new_n711), .B2(new_n636), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n683), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n680), .B1(new_n714), .B2(G1), .ZN(G364));
  INV_X1    g0515(.A(new_n677), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n261), .A2(G20), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n203), .B1(new_n717), .B2(G45), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n663), .A2(G330), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n665), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT92), .Z(new_n723));
  NOR2_X1   g0523(.A1(new_n676), .A2(new_n275), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G355), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G116), .B2(new_n207), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n676), .A2(new_n512), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n225), .B2(new_n288), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n246), .A2(G45), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT93), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n226), .B1(G20), .B2(new_n498), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n720), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n734), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n663), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n204), .A2(new_n308), .A3(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n579), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n383), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n743), .A2(G58), .B1(G77), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n204), .A2(new_n308), .A3(new_n337), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n747), .A2(KEYINPUT95), .A3(new_n383), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT95), .B1(new_n747), .B2(new_n383), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n746), .A2(KEYINPUT94), .B1(new_n751), .B2(G68), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(KEYINPUT94), .B2(new_n746), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n579), .A2(new_n747), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n275), .B1(new_n755), .B2(G50), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n204), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n383), .A3(new_n337), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G159), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT32), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n383), .A2(G179), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n204), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n757), .A2(new_n383), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n764), .A2(G97), .B1(new_n766), .B2(G107), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n213), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n760), .B2(KEYINPUT32), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n756), .A2(new_n761), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n754), .B(KEYINPUT96), .Z(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n773), .B1(new_n750), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n744), .A2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n512), .B(new_n777), .C1(G329), .C2(new_n759), .ZN(new_n778));
  INV_X1    g0578(.A(new_n768), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n764), .A2(G294), .B1(new_n779), .B2(G303), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n743), .A2(G322), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(G283), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n778), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n753), .A2(new_n771), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n738), .B(new_n740), .C1(new_n735), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n723), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n335), .A2(new_n660), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n320), .A2(new_n334), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n330), .B(new_n331), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n660), .B1(new_n790), .B2(new_n323), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n789), .B1(new_n791), .B2(new_n339), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n681), .B(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n720), .B1(new_n795), .B2(new_n708), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n708), .B2(new_n795), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n735), .A2(new_n732), .ZN(new_n798));
  INV_X1    g0598(.A(G132), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n512), .B1(new_n758), .B2(new_n799), .C1(new_n211), .C2(new_n765), .ZN(new_n800));
  INV_X1    g0600(.A(G58), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n763), .A2(new_n801), .B1(new_n768), .B2(new_n250), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n755), .A2(G137), .B1(new_n745), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(G143), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n742), .C1(new_n750), .C2(new_n248), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n800), .B(new_n802), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n755), .A2(G303), .B1(new_n745), .B2(G116), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n750), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT97), .Z(new_n812));
  OAI22_X1  g0612(.A1(new_n213), .A2(new_n765), .B1(new_n768), .B2(new_n520), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n275), .B1(new_n758), .B2(new_n776), .C1(new_n763), .C2(new_n562), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(G294), .C2(new_n743), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n807), .A2(new_n808), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n735), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n720), .B1(G77), .B2(new_n798), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT98), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n733), .B2(new_n794), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n797), .A2(new_n820), .ZN(G384));
  INV_X1    g0621(.A(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n611), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n823), .A2(G20), .A3(G116), .A4(new_n227), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT99), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n825), .B1(new_n822), .B2(new_n611), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT36), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n225), .B(G77), .C1(new_n801), .C2(new_n211), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n250), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n203), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n717), .A2(new_n203), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n412), .A2(new_n415), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT16), .B1(new_n834), .B2(new_n420), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n447), .B1(new_n835), .B2(new_n417), .ZN(new_n836));
  INV_X1    g0636(.A(new_n657), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n459), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n445), .A2(new_n836), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n450), .A2(new_n837), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n459), .C1(new_n426), .C2(new_n443), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(KEYINPUT37), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  INV_X1    g0645(.A(new_n838), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n464), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n845), .B1(new_n464), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT38), .B(new_n844), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(KEYINPUT102), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n854), .A3(new_n850), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n464), .A2(new_n450), .A3(new_n837), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n843), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n850), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n394), .A2(new_n659), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT100), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n356), .A2(new_n866), .A3(new_n659), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n356), .B2(new_n659), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n387), .B2(new_n394), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n387), .A2(new_n394), .A3(new_n869), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n630), .B1(new_n634), .B2(new_n635), .C1(new_n644), .C2(KEYINPUT88), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n641), .A2(new_n644), .A3(KEYINPUT88), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n660), .B(new_n794), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(new_n788), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n853), .A3(new_n855), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n651), .A2(new_n657), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n865), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n465), .B1(new_n683), .B2(new_n713), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n652), .A2(new_n310), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n882), .B(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n387), .A2(new_n869), .A3(new_n394), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n870), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n794), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n627), .A2(KEYINPUT31), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n694), .A2(new_n659), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n702), .A2(new_n703), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n853), .A2(new_n855), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n852), .B2(new_n860), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n896), .A2(new_n897), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n892), .A2(new_n894), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n900), .A2(new_n629), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  INV_X1    g0703(.A(G330), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n833), .B1(new_n886), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT103), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n906), .A2(new_n907), .B1(new_n886), .B2(new_n905), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n832), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT104), .ZN(G367));
  OAI21_X1  g0711(.A(new_n736), .B1(new_n728), .B2(new_n238), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n676), .B2(new_n326), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n719), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n505), .A2(new_n660), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(new_n630), .A3(new_n631), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n630), .B2(new_n916), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n772), .A2(new_n776), .ZN(new_n919));
  INV_X1    g0719(.A(G317), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n275), .B1(new_n758), .B2(new_n920), .C1(new_n744), .C2(new_n810), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n779), .A2(KEYINPUT46), .A3(G116), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT46), .B1(new_n779), .B2(G116), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n751), .A2(G294), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n765), .A2(new_n562), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n763), .A2(new_n520), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n743), .C2(G303), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n919), .A2(new_n924), .A3(new_n925), .A4(new_n928), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n742), .A2(new_n248), .B1(new_n321), .B2(new_n765), .ZN(new_n930));
  INV_X1    g0730(.A(G137), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n512), .B1(new_n758), .B2(new_n931), .C1(new_n744), .C2(new_n250), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n763), .A2(new_n211), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n768), .A2(new_n801), .ZN(new_n934));
  NOR4_X1   g0734(.A1(new_n930), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n935), .B1(new_n804), .B2(new_n772), .C1(new_n400), .C2(new_n750), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT47), .Z(new_n938));
  OAI221_X1 g0738(.A(new_n914), .B1(new_n739), .B2(new_n918), .C1(new_n938), .C2(new_n817), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n718), .B(KEYINPUT108), .ZN(new_n940));
  MUX2_X1   g0740(.A(new_n557), .B(new_n668), .S(new_n670), .Z(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(new_n664), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n714), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n617), .A2(new_n659), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n622), .A2(new_n624), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(new_n624), .C2(new_n660), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n672), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT44), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n672), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT106), .Z(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(KEYINPUT45), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n669), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT107), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n943), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n953), .B2(new_n954), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n714), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n677), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n940), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n946), .A2(new_n947), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n624), .B1(new_n965), .B2(new_n556), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n948), .A2(new_n671), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n966), .A2(new_n660), .B1(new_n967), .B2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(KEYINPUT42), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n956), .A2(new_n948), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n939), .B1(new_n964), .B2(new_n976), .ZN(G387));
  NOR2_X1   g0777(.A1(new_n714), .A2(new_n942), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n943), .A2(new_n978), .A3(new_n716), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n668), .A2(new_n739), .ZN(new_n980));
  INV_X1    g0780(.A(new_n675), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n252), .A2(G50), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g0784(.A(G45), .B1(G68), .B2(G77), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT111), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n984), .B(new_n985), .C1(new_n675), .C2(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n727), .B1(new_n235), .B2(new_n288), .C1(new_n982), .C2(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n675), .A2(new_n724), .B1(new_n520), .B2(new_n676), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT110), .Z(new_n990));
  AOI21_X1  g0790(.A(new_n737), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n980), .A2(new_n719), .A3(new_n991), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n275), .B(new_n926), .C1(G150), .C2(new_n759), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G50), .A2(new_n743), .B1(new_n755), .B2(G159), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n745), .A2(G68), .B1(new_n779), .B2(G77), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n326), .A2(new_n764), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n253), .B2(new_n751), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT112), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n512), .B1(new_n759), .B2(G326), .ZN(new_n1000));
  INV_X1    g0800(.A(G294), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n763), .A2(new_n810), .B1(new_n768), .B2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n743), .A2(G317), .B1(G303), .B2(new_n745), .ZN(new_n1003));
  INV_X1    g0803(.A(G322), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n776), .B2(new_n750), .C1(new_n772), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT48), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1000), .B1(new_n559), .B2(new_n765), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n999), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n992), .B1(new_n735), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n942), .A2(new_n940), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT109), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n979), .A2(new_n1013), .A3(new_n1015), .ZN(G393));
  XNOR2_X1  g0816(.A(new_n955), .B(new_n669), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n940), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n243), .A2(new_n727), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n736), .B1(new_n562), .B2(new_n207), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n720), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n512), .B1(new_n758), .B2(new_n804), .C1(new_n213), .C2(new_n765), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n763), .A2(new_n321), .B1(new_n768), .B2(new_n211), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n253), .C2(new_n745), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n250), .B2(new_n750), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n248), .A2(new_n754), .B1(new_n742), .B2(new_n400), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT51), .Z(new_n1027));
  OAI22_X1  g0827(.A1(new_n763), .A2(new_n559), .B1(new_n768), .B2(new_n810), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n275), .B1(new_n758), .B2(new_n1004), .C1(new_n520), .C2(new_n765), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G294), .C2(new_n745), .ZN(new_n1030));
  INV_X1    g0830(.A(G303), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(new_n1031), .B2(new_n750), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n776), .A2(new_n742), .B1(new_n754), .B2(new_n920), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT52), .Z(new_n1034));
  OAI22_X1  g0834(.A1(new_n1025), .A2(new_n1027), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT113), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n1021), .B1(new_n1036), .B2(new_n735), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n948), .B2(new_n739), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1017), .A2(new_n943), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n677), .B1(new_n959), .B2(new_n960), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1018), .B(new_n1038), .C1(new_n1039), .C2(new_n1040), .ZN(G390));
  NAND3_X1  g0841(.A1(new_n900), .A2(G330), .A3(new_n629), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1043), .A2(new_n883), .A3(new_n884), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n788), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n681), .B2(new_n794), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n887), .A2(new_n870), .A3(new_n793), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(G330), .C1(new_n695), .C2(new_n893), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(G330), .B(new_n794), .C1(new_n695), .C2(new_n707), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n873), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1049), .B1(new_n1051), .B2(KEYINPUT115), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT115), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1053), .A3(new_n873), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1046), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1050), .A2(new_n873), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n792), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n712), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n1045), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n873), .B(KEYINPUT114), .ZN(new_n1060));
  OAI211_X1 g0860(.A(G330), .B(new_n794), .C1(new_n695), .C2(new_n893), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1056), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1044), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n864), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1046), .B2(new_n873), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n856), .A2(new_n1066), .A3(new_n862), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n861), .C1(new_n1060), .C2(new_n1059), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n1067), .A2(new_n1056), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1048), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1049), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1056), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1050), .A2(new_n1053), .A3(new_n873), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1053), .B1(new_n1050), .B2(new_n873), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1075), .A2(new_n1076), .A3(new_n1049), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1077), .B2(new_n1046), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1067), .A2(new_n1068), .A3(new_n1056), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n1078), .A3(new_n1079), .A4(new_n1044), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1071), .A2(new_n1080), .A3(new_n677), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n720), .B1(new_n798), .B2(new_n253), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT54), .B(G143), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n751), .A2(G137), .B1(new_n745), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT117), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT117), .ZN(new_n1087));
  INV_X1    g0887(.A(G128), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1088), .A2(new_n754), .B1(new_n742), .B2(new_n799), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n275), .B1(new_n759), .B2(G125), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n250), .B2(new_n765), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(G159), .C2(new_n764), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n768), .A2(new_n248), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT53), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1086), .A2(new_n1087), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n755), .A2(G283), .B1(new_n745), .B2(G97), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n520), .B2(new_n750), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT118), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n765), .A2(new_n211), .B1(new_n758), .B2(new_n1001), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n742), .A2(new_n559), .B1(new_n321), .B2(new_n763), .ZN(new_n1101));
  OR4_X1    g0901(.A1(new_n512), .A2(new_n1100), .A3(new_n769), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1095), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1082), .B1(new_n1103), .B2(new_n735), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n863), .B2(new_n733), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n940), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(KEYINPUT116), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(KEYINPUT116), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1081), .B(new_n1105), .C1(new_n1108), .C2(new_n1109), .ZN(G378));
  INV_X1    g0910(.A(KEYINPUT57), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n896), .A2(new_n897), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n904), .B1(new_n895), .B2(new_n898), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n307), .A2(new_n310), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n268), .A2(new_n837), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1117), .B(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1112), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n882), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n880), .B1(new_n864), .B2(new_n863), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1112), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1120), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1044), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1106), .B2(new_n1078), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1111), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1080), .A2(new_n1044), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT121), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1124), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n882), .A2(new_n1122), .A3(new_n1123), .A4(KEYINPUT121), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n1135), .A3(KEYINPUT57), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1137), .A3(new_n677), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1121), .A2(new_n733), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n720), .B1(new_n798), .B2(G50), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n512), .A2(G41), .ZN(new_n1141));
  AOI211_X1 g0941(.A(G50), .B(new_n1141), .C1(new_n254), .C2(new_n287), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n765), .A2(new_n801), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n742), .A2(new_n520), .B1(new_n321), .B2(new_n768), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G116), .C2(new_n755), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1141), .B1(new_n810), .B2(new_n758), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n933), .B(new_n1146), .C1(new_n326), .C2(new_n745), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(new_n562), .C2(new_n750), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT58), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G33), .B(G41), .C1(new_n759), .C2(G124), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n768), .A2(new_n1083), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT120), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n755), .A2(G125), .B1(G150), .B2(new_n764), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n1088), .B2(new_n742), .C1(new_n931), .C2(new_n744), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(G132), .C2(new_n751), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT59), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1151), .B1(new_n400), .B2(new_n765), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1150), .B1(new_n1149), .B2(new_n1148), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1140), .B1(new_n1160), .B2(new_n735), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1139), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n940), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1138), .A2(new_n1165), .ZN(G375));
  NAND2_X1  g0966(.A1(new_n1060), .A2(new_n732), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n720), .B1(new_n798), .B2(G68), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n742), .A2(new_n931), .B1(new_n400), .B2(new_n768), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G150), .B2(new_n745), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n751), .A2(new_n1084), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n275), .B(new_n1143), .C1(G128), .C2(new_n759), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n755), .A2(G132), .B1(G50), .B2(new_n764), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n754), .A2(new_n1001), .B1(new_n520), .B2(new_n744), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G283), .B2(new_n743), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n751), .A2(G116), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n512), .B1(new_n766), .B2(G77), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n996), .A4(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n758), .A2(new_n1031), .B1(new_n768), .B2(new_n562), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT122), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1174), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1168), .B1(new_n1182), .B2(new_n735), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1078), .A2(new_n940), .B1(new_n1167), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1064), .A2(new_n963), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1055), .A2(new_n1063), .A3(new_n1044), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(G381));
  INV_X1    g0987(.A(G390), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n964), .A2(new_n976), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n939), .A4(new_n1190), .ZN(new_n1191));
  OR4_X1    g0991(.A1(G378), .A2(new_n1191), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g0992(.A1(new_n658), .A2(G213), .ZN(new_n1193));
  OR3_X1    g0993(.A1(G375), .A2(G378), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(G407), .A2(G213), .A3(new_n1194), .ZN(G409));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1164), .A2(new_n963), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n1131), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n962), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1133), .A3(KEYINPUT123), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1163), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT124), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1135), .A2(new_n1202), .A3(new_n1136), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n940), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G378), .B1(new_n1201), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1138), .A2(G378), .A3(new_n1165), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1193), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n658), .A2(G213), .A3(G2897), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1046), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1214), .A2(new_n1130), .A3(KEYINPUT60), .A4(new_n1074), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1078), .B2(new_n1044), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n677), .B(new_n1215), .C1(new_n1218), .C2(new_n1186), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1219), .A2(G384), .A3(new_n1184), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G384), .B1(new_n1219), .B2(new_n1184), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1211), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT127), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(KEYINPUT127), .B(new_n1211), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1186), .B1(new_n1064), .B2(new_n1216), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n677), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1184), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1219), .A2(G384), .A3(new_n1184), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1210), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1230), .A2(KEYINPUT126), .A3(new_n1231), .A4(new_n1210), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1224), .A2(new_n1225), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT61), .B1(new_n1209), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(G378), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1200), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT123), .B1(new_n1199), .B2(new_n1133), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1162), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1205), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n940), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1242), .A2(new_n1203), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1238), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1138), .A2(G378), .A3(new_n1165), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1193), .A4(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1193), .B(new_n1249), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1237), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1189), .A2(G390), .A3(new_n939), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1188), .A2(G387), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(G393), .B(new_n786), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1253), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1251), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1193), .A4(new_n1249), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1261), .A2(new_n1237), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(G405));
  XNOR2_X1  g1068(.A(G375), .B(G378), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1249), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1262), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(new_n1261), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G402));
endmodule


