//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT82), .Z(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT77), .B1(new_n205), .B2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT76), .B1(new_n207), .B2(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(new_n207), .A3(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(new_n205), .A3(G148gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n206), .A2(new_n208), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT2), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n207), .A2(G141gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n205), .A2(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n215), .A2(new_n214), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n213), .A2(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G197gat), .B(G204gat), .Z(new_n223));
  AOI21_X1  g022(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT83), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n231), .B(new_n232), .C1(KEYINPUT83), .C2(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n222), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(new_n234), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n229), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n204), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n229), .B2(new_n232), .ZN(new_n239));
  OAI211_X1 g038(.A(G228gat), .B(G233gat), .C1(new_n239), .C2(new_n222), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G78gat), .B(G106gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G22gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT31), .B(G50gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n241), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT67), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  OR3_X1    g053(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n254), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT23), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(G169gat), .B2(G176gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n266), .A3(new_n257), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n248), .A3(KEYINPUT64), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(G183gat), .B2(G190gat), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n267), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT65), .B1(new_n277), .B2(KEYINPUT25), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n264), .A2(new_n266), .A3(new_n257), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n252), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(new_n269), .A3(new_n271), .A4(new_n273), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n274), .A2(new_n275), .A3(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n289), .A2(new_n267), .A3(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n261), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g091(.A(KEYINPUT66), .B(new_n290), .C1(new_n278), .C2(new_n286), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n260), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295));
  INV_X1    g094(.A(G113gat), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g098(.A1(G113gat), .A2(G120gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n303));
  INV_X1    g102(.A(G127gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(G134gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n302), .B1(new_n301), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n295), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(G113gat), .B2(G120gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n300), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(KEYINPUT71), .A3(new_n306), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n294), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G227gat), .ZN(new_n320));
  INV_X1    g119(.A(G233gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n323));
  AOI211_X1 g122(.A(KEYINPUT65), .B(KEYINPUT25), .C1(new_n279), .C2(new_n282), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n291), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n287), .A2(new_n261), .A3(new_n291), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n316), .A4(new_n260), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n319), .A2(new_n322), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G15gat), .B(G43gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n330), .B(KEYINPUT32), .C1(new_n332), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n329), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n320), .B2(new_n321), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT34), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT34), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n344), .C1(new_n320), .C2(new_n321), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n337), .A2(new_n343), .A3(new_n345), .A4(new_n339), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n337), .A2(new_n339), .B1(new_n343), .B2(new_n345), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n246), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n309), .A2(new_n222), .A3(new_n315), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n307), .A2(new_n308), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n213), .A2(new_n216), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n220), .A2(new_n221), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  OAI22_X1  g161(.A1(new_n355), .A2(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n357), .A3(new_n236), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n363), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n365), .A2(new_n366), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n371), .A3(new_n356), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n361), .A2(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n355), .B2(new_n356), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n360), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n222), .B1(new_n307), .B2(new_n308), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT80), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n380), .A3(new_n360), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n367), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n382), .A2(KEYINPUT5), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n369), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385));
  INV_X1    g184(.A(G85gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT0), .B(G57gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n354), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT6), .B1(new_n384), .B2(new_n390), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n355), .A2(new_n356), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT79), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n373), .A3(new_n372), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n396), .B2(new_n370), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT81), .B(new_n389), .C1(new_n397), .C2(new_n369), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n391), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT6), .B(new_n389), .C1(new_n397), .C2(new_n369), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n325), .A2(new_n260), .ZN(new_n402));
  AND2_X1   g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n260), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n326), .B2(new_n327), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n403), .A2(KEYINPUT29), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n404), .B(new_n230), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT74), .B(G64gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n325), .A2(new_n260), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n406), .A2(new_n403), .B1(new_n415), .B2(new_n407), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n409), .B(new_n414), .C1(new_n416), .C2(new_n230), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n328), .A2(new_n260), .A3(new_n403), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n402), .A2(new_n408), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n229), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n418), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(KEYINPUT30), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n401), .A2(new_n420), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n202), .B1(new_n353), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(KEYINPUT30), .ZN(new_n430));
  INV_X1    g229(.A(new_n424), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n420), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n426), .B2(new_n420), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n348), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n437), .A2(new_n246), .A3(new_n350), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n389), .B1(new_n397), .B2(new_n369), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n392), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT35), .B1(new_n440), .B2(new_n400), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n436), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT36), .B1(new_n347), .B2(new_n348), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n349), .A2(new_n352), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(KEYINPUT36), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n246), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n367), .B1(new_n379), .B2(new_n381), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n363), .A2(new_n365), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n367), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n448), .A3(new_n367), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n390), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n447), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n454), .A2(KEYINPUT40), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n439), .B1(new_n454), .B2(KEYINPUT40), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n426), .A2(new_n434), .A3(new_n420), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n440), .A2(new_n400), .A3(new_n417), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT86), .A3(new_n229), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n416), .A2(new_n230), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT86), .B1(new_n462), .B2(new_n229), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n409), .B(new_n468), .C1(new_n416), .C2(new_n230), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n414), .A2(KEYINPUT38), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n413), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n423), .B2(new_n409), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT38), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n461), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n246), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n446), .B1(new_n460), .B2(new_n478), .ZN(new_n479));
  OAI22_X1  g278(.A1(new_n429), .A2(new_n442), .B1(new_n445), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT91), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(G1gat), .ZN(new_n484));
  INV_X1    g283(.A(G8gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n481), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G1gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n484), .B2(new_n489), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G71gat), .B(G78gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(KEYINPUT94), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(G57gat), .B(G64gat), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(KEYINPUT94), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT94), .B(new_n493), .C1(new_n496), .C2(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n492), .B1(new_n504), .B2(new_n502), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G231gat), .A2(G233gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(new_n268), .ZN(new_n508));
  INV_X1    g307(.A(G211gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n506), .A2(new_n510), .ZN(new_n512));
  XOR2_X1   g311(.A(G127gat), .B(G155gat), .Z(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n511), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n511), .B2(new_n512), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT41), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT95), .ZN(new_n523));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  INV_X1    g326(.A(G92gat), .ZN(new_n528));
  AOI22_X1  g327(.A1(KEYINPUT8), .A2(new_n527), .B1(new_n386), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n386), .B2(new_n528), .ZN(new_n531));
  NAND3_X1  g330(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G99gat), .B(G106gat), .Z(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT96), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT90), .B(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT14), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n544), .B1(KEYINPUT89), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(KEYINPUT89), .B2(new_n547), .ZN(new_n549));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n547), .A2(new_n551), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  INV_X1    g353(.A(new_n550), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n544), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n549), .A2(new_n552), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(KEYINPUT41), .B2(new_n521), .ZN(new_n559));
  XOR2_X1   g358(.A(G190gat), .B(G218gat), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n541), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n561), .B1(new_n559), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n526), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(new_n525), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT97), .B1(new_n520), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n519), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT10), .B(new_n501), .C1(new_n538), .C2(new_n540), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n501), .A2(new_n537), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n499), .B(new_n500), .C1(new_n536), .C2(new_n535), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT10), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n577), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT98), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n585));
  AOI211_X1 g384(.A(new_n585), .B(new_n577), .C1(new_n578), .C2(new_n582), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n579), .A2(new_n580), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(new_n577), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  INV_X1    g394(.A(new_n583), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n577), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n573), .A2(new_n575), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n573), .A2(KEYINPUT99), .A3(new_n575), .A4(new_n599), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n549), .A2(new_n552), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n556), .A2(new_n553), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n605), .A2(new_n606), .B1(new_n490), .B2(new_n491), .ZN(new_n607));
  INV_X1    g406(.A(new_n491), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n557), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n604), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n608), .B(new_n609), .C1(new_n557), .C2(KEYINPUT17), .ZN(new_n617));
  INV_X1    g416(.A(new_n563), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n612), .B(new_n607), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT18), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n562), .A2(new_n492), .A3(new_n563), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n612), .A4(new_n607), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n611), .A2(new_n604), .A3(new_n614), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n616), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n205), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT88), .B(G113gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n635));
  AOI211_X1 g434(.A(KEYINPUT92), .B(new_n613), .C1(new_n607), .C2(new_n610), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n615), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n637), .A2(new_n623), .A3(new_n621), .A4(new_n632), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n625), .A2(KEYINPUT93), .A3(new_n633), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n480), .A2(new_n602), .A3(new_n603), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n401), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n488), .ZN(G1324gat));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  INV_X1    g444(.A(new_n436), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT16), .B(G8gat), .Z(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT42), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n646), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(G8gat), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n648), .B2(new_n652), .ZN(G1325gat));
  NOR2_X1   g452(.A1(new_n437), .A2(new_n350), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G15gat), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT100), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  INV_X1    g457(.A(new_n445), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n642), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n477), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n480), .A2(new_n572), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n436), .A2(new_n438), .A3(new_n441), .ZN(new_n669));
  AOI211_X1 g468(.A(new_n427), .B(new_n246), .C1(new_n349), .C2(new_n352), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n202), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n455), .A2(new_n456), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n433), .B2(new_n435), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n423), .A2(new_n409), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT37), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n413), .A3(new_n469), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n676), .A2(KEYINPUT38), .B1(new_n467), .B2(new_n471), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n246), .B1(new_n677), .B2(new_n461), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT36), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n349), .B2(new_n352), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n679), .B(new_n446), .C1(new_n681), .C2(new_n443), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n571), .B1(new_n671), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n639), .A2(new_n640), .ZN(new_n687));
  INV_X1    g486(.A(new_n599), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n519), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n401), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(new_n542), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n683), .A2(new_n689), .ZN(new_n693));
  INV_X1    g492(.A(new_n401), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n542), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT102), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n692), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n693), .A2(new_n543), .A3(new_n646), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT46), .Z(new_n703));
  OAI21_X1  g502(.A(G36gat), .B1(new_n690), .B2(new_n436), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1329gat));
  OAI21_X1  g504(.A(G43gat), .B1(new_n690), .B2(new_n659), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n693), .A2(new_n711), .A3(new_n654), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n706), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n706), .B2(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n712), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT104), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n718), .A2(new_n708), .A3(new_n707), .A4(new_n713), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1330gat));
  OAI21_X1  g519(.A(G50gat), .B1(new_n690), .B2(new_n477), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT48), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G50gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n693), .A2(new_n724), .A3(new_n246), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n723), .B(new_n726), .ZN(G1331gat));
  NAND3_X1  g526(.A1(new_n573), .A2(new_n575), .A3(new_n687), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n599), .B(new_n728), .C1(new_n671), .C2(new_n682), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n694), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n646), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n654), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT106), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(KEYINPUT106), .ZN(new_n738));
  AOI21_X1  g537(.A(G71gat), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n729), .A2(new_n445), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(G71gat), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n729), .A2(new_n246), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT107), .B(G78gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n687), .A2(new_n520), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT108), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n599), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n686), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n401), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT51), .B1(new_n683), .B2(new_n747), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n480), .A2(KEYINPUT51), .A3(new_n572), .A4(new_n747), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n683), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n747), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n688), .A2(new_n694), .A3(new_n386), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n751), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  NOR3_X1   g561(.A1(new_n436), .A2(G92gat), .A3(new_n599), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n686), .A2(new_n646), .A3(new_n749), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n752), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n758), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n770), .A2(new_n763), .B1(new_n765), .B2(G92gat), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n764), .A2(new_n768), .B1(new_n767), .B2(new_n771), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n750), .B2(new_n659), .ZN(new_n773));
  INV_X1    g572(.A(G99gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n654), .A2(new_n774), .A3(new_n688), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n760), .B2(new_n775), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g576(.A(G106gat), .B1(new_n750), .B2(new_n477), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n477), .A2(new_n599), .A3(G106gat), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n777), .B(new_n778), .C1(new_n760), .C2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n770), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT111), .B1(new_n784), .B2(new_n780), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n778), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT53), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n786), .B2(KEYINPUT53), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n781), .B1(new_n788), .B2(new_n789), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n578), .A2(new_n582), .A3(new_n577), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(KEYINPUT54), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n584), .B2(new_n586), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n595), .B1(new_n583), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n593), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n795), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n797), .A2(KEYINPUT113), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n593), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n800), .A2(new_n640), .A3(new_n639), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n612), .B1(new_n622), .B2(new_n607), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n611), .A2(new_n614), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n631), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n638), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n599), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n572), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n800), .A2(new_n802), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(new_n571), .A3(new_n807), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n520), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n728), .A2(new_n688), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n646), .A2(new_n401), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n353), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n296), .A3(new_n641), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n438), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n687), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1340gat));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n297), .A3(new_n688), .ZN(new_n823));
  OAI21_X1  g622(.A(G120gat), .B1(new_n820), .B2(new_n599), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1341gat));
  AOI21_X1  g624(.A(G127gat), .B1(new_n818), .B2(new_n519), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n820), .A2(new_n304), .A3(new_n520), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(G1342gat));
  INV_X1    g627(.A(G134gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n829), .A3(new_n572), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n817), .A2(new_n438), .A3(new_n572), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n832), .B(new_n833), .C1(new_n829), .C2(new_n834), .ZN(G1343gat));
  NAND2_X1  g634(.A1(new_n659), .A2(new_n815), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n477), .B1(new_n812), .B2(new_n813), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n799), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT115), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n798), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n797), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n841), .A2(KEYINPUT116), .A3(new_n798), .A4(new_n842), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n641), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n572), .B1(new_n848), .B2(new_n808), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n520), .B1(new_n849), .B2(new_n811), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n477), .B1(new_n850), .B2(new_n813), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n839), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G141gat), .B1(new_n852), .B2(new_n687), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n659), .A2(new_n246), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n816), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n205), .A3(new_n641), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n853), .A2(new_n861), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n862), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n860), .B1(new_n864), .B2(new_n854), .ZN(G1344gat));
  INV_X1    g664(.A(new_n852), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n207), .C1(new_n866), .C2(new_n688), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n602), .A2(new_n603), .A3(new_n687), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n477), .B1(new_n850), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n838), .B(new_n477), .C1(new_n812), .C2(new_n813), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n814), .A2(new_n246), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT119), .B1(new_n874), .B2(new_n838), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n836), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(G148gat), .A3(new_n688), .A4(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n856), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n207), .B1(new_n879), .B2(new_n599), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n867), .B1(new_n881), .B2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g681(.A(G155gat), .B1(new_n856), .B2(new_n519), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n519), .A2(G155gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n866), .B2(new_n884), .ZN(G1346gat));
  NOR4_X1   g684(.A1(new_n816), .A2(G162gat), .A3(new_n571), .A4(new_n855), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT120), .Z(new_n887));
  OAI21_X1  g686(.A(G162gat), .B1(new_n852), .B2(new_n571), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1347gat));
  AOI211_X1 g688(.A(new_n694), .B(new_n436), .C1(new_n812), .C2(new_n813), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n353), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n262), .A3(new_n641), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n438), .ZN(new_n893));
  OAI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n687), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1348gat));
  NOR3_X1   g694(.A1(new_n893), .A2(new_n263), .A3(new_n599), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n891), .A2(new_n688), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n263), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(KEYINPUT121), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(KEYINPUT121), .B2(new_n899), .ZN(G1349gat));
  NAND3_X1  g700(.A1(new_n891), .A2(new_n247), .A3(new_n519), .ZN(new_n902));
  OAI21_X1  g701(.A(G183gat), .B1(new_n893), .B2(new_n520), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n904), .B(new_n905), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n893), .B2(new_n571), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT61), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n248), .A3(new_n572), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1351gat));
  OAI22_X1  g709(.A1(new_n871), .A2(new_n872), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n838), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT124), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n870), .A2(new_n875), .A3(new_n873), .A4(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n445), .A2(new_n694), .A3(new_n436), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n687), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n837), .A2(new_n916), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n687), .A2(G197gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1352gat));
  NAND4_X1  g720(.A1(new_n913), .A2(new_n915), .A3(new_n688), .A4(new_n916), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT125), .B(G204gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n919), .A2(new_n599), .A3(new_n923), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n519), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n509), .B1(new_n876), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT63), .ZN(new_n935));
  INV_X1    g734(.A(new_n919), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n509), .A3(new_n519), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1354gat));
  NAND2_X1  g737(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n913), .A2(new_n915), .A3(new_n940), .A4(new_n916), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n572), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G218gat), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n919), .A2(G218gat), .A3(new_n571), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


