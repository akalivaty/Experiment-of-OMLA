//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1339,
    new_n1340, new_n1341, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1419,
    new_n1420, new_n1421, new_n1422;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND3_X1  g0015(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  INV_X1    g0045(.A(G45), .ZN(new_n246));
  AOI21_X1  g0046(.A(G1), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  AND3_X1   g0049(.A1(new_n247), .A2(new_n249), .A3(G274), .ZN(new_n250));
  INV_X1    g0050(.A(new_n249), .ZN(new_n251));
  INV_X1    g0051(.A(G226), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n251), .A2(new_n247), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n257), .A3(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(G1698), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n258), .B1(new_n206), .B2(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI211_X1 g0061(.A(new_n250), .B(new_n253), .C1(new_n261), .C2(new_n251), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G190), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n209), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n269), .A2(new_n272), .B1(new_n273), .B2(new_n265), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(new_n210), .A3(new_n279), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n278), .A2(new_n280), .B1(new_n284), .B2(G150), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n205), .B2(new_n210), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n275), .B1(new_n286), .B2(new_n268), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n263), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G200), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n262), .A2(new_n291), .B1(new_n287), .B2(KEYINPUT9), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n288), .B1(new_n262), .B2(G169), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n262), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n268), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n284), .A2(G50), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n280), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n307), .A2(KEYINPUT11), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(KEYINPUT11), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n310), .A2(new_n311), .B1(new_n269), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G33), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n316), .A2(new_n318), .A3(G232), .A4(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  OR2_X1    g0120(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n321), .A2(new_n316), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n319), .B(new_n320), .C1(new_n323), .C2(new_n252), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n251), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n247), .A2(new_n249), .A3(G274), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n249), .A2(G238), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n315), .B1(new_n335), .B2(G169), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n325), .B2(new_n330), .ZN(new_n337));
  AOI211_X1 g0137(.A(KEYINPUT13), .B(new_n329), .C1(new_n324), .C2(new_n251), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n315), .B(G169), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(G179), .A3(new_n334), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n314), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n332), .A2(G190), .A3(new_n334), .ZN(new_n344));
  INV_X1    g0144(.A(new_n314), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n337), .A2(new_n338), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n291), .ZN(new_n349));
  OAI211_X1 g0149(.A(KEYINPUT71), .B(G200), .C1(new_n337), .C2(new_n338), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n278), .A2(new_n270), .ZN(new_n354));
  INV_X1    g0154(.A(new_n278), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n354), .A2(new_n269), .B1(new_n265), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT72), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(G58), .A3(G68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n360), .A3(new_n203), .ZN(new_n361));
  AOI22_X1  g0161(.A1(G20), .A2(new_n361), .B1(new_n284), .B2(G159), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n317), .A2(G33), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n210), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n316), .A2(new_n318), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(G20), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n362), .C1(new_n369), .C2(new_n202), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n268), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n316), .A2(new_n318), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n368), .B1(new_n316), .B2(new_n372), .ZN(new_n374));
  AOI21_X1  g0174(.A(G20), .B1(new_n316), .B2(new_n318), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n373), .A2(new_n374), .B1(new_n375), .B2(KEYINPUT7), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G68), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT16), .B1(new_n377), .B2(new_n362), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n356), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n323), .A2(new_n259), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n316), .A2(new_n318), .A3(G226), .A4(G1698), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n251), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n249), .A2(G232), .A3(new_n327), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n249), .A2(new_n327), .A3(KEYINPUT74), .A4(G232), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n250), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(G200), .B1(new_n384), .B2(new_n389), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n353), .B1(new_n379), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n384), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n291), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(G190), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n316), .A2(new_n318), .A3(new_n372), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n368), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n366), .B1(new_n257), .B2(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n202), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n361), .A2(G20), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n284), .A2(G159), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n268), .A3(new_n370), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n408), .A4(new_n356), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n394), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n387), .A2(new_n388), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n326), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n381), .A2(new_n382), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n256), .A2(new_n257), .A3(G223), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n249), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G169), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n384), .A2(new_n389), .A3(G179), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n379), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT18), .B1(new_n379), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n284), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n355), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  INV_X1    g0226(.A(new_n280), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n210), .B2(new_n206), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n268), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n270), .A2(G77), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n269), .A2(new_n431), .B1(new_n206), .B2(new_n265), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n256), .A2(new_n257), .A3(G232), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n435), .B1(new_n436), .B2(new_n257), .C1(new_n219), .C2(new_n260), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n251), .ZN(new_n438));
  INV_X1    g0238(.A(G244), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n251), .A2(new_n247), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n250), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(KEYINPUT69), .B(new_n434), .C1(new_n442), .C2(new_n291), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT69), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n291), .B1(new_n438), .B2(new_n441), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n433), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n441), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n443), .B(new_n446), .C1(new_n390), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G169), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n434), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT70), .B1(new_n442), .B2(new_n298), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT70), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n447), .A2(new_n452), .A3(G179), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n303), .A2(new_n352), .A3(new_n423), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(G303), .B1(new_n363), .B2(new_n364), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n316), .A2(new_n318), .A3(G264), .A4(G1698), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n256), .A2(new_n257), .A3(G257), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT80), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(KEYINPUT80), .A3(new_n459), .A4(new_n458), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n251), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n246), .A2(G1), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G270), .A3(new_n249), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(G274), .A3(new_n249), .A4(new_n467), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n465), .A2(new_n466), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n458), .B(new_n459), .C1(new_n323), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n249), .B1(new_n480), .B2(new_n463), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT81), .B1(new_n481), .B2(new_n474), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n210), .C1(G33), .C2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(new_n268), .C1(new_n210), .C2(G116), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT20), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n264), .A2(G116), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n269), .B1(G1), .B2(new_n279), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n484), .A2(KEYINPUT82), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT82), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n291), .B1(new_n476), .B2(new_n482), .ZN(new_n498));
  INV_X1    g0298(.A(new_n495), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n476), .A2(new_n482), .A3(G190), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  INV_X1    g0303(.A(new_n492), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G107), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n264), .A2(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT25), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n436), .A3(G20), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT24), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n509), .A2(new_n511), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n316), .A2(new_n318), .A3(new_n210), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n257), .A2(new_n518), .A3(new_n210), .A4(G87), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n513), .A2(KEYINPUT24), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n520), .B(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n508), .B1(new_n522), .B2(new_n268), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n321), .A2(G250), .A3(new_n322), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G257), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n367), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G294), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n279), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n251), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n470), .A2(new_n249), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G264), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n531), .A3(new_n473), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n449), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n529), .A2(new_n531), .A3(new_n298), .A4(new_n473), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n503), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n517), .A2(new_n519), .ZN(new_n538));
  INV_X1    g0338(.A(new_n515), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n521), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n521), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n541), .B(new_n515), .C1(new_n517), .C2(new_n519), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n268), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n505), .A3(new_n507), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n544), .A3(KEYINPUT84), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n532), .A2(new_n291), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n529), .A2(new_n531), .A3(new_n390), .A4(new_n473), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(KEYINPUT85), .A3(new_n547), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n547), .A2(KEYINPUT85), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n523), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n536), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n471), .A2(G179), .A3(new_n473), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n499), .A2(new_n465), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(G169), .B1(new_n489), .B2(new_n494), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n466), .B1(new_n465), .B2(new_n475), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n481), .A2(KEYINPUT81), .A3(new_n474), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n483), .A2(new_n561), .A3(new_n556), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n554), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n502), .A2(new_n551), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT4), .A4(G244), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n565), .A2(new_n485), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n323), .B2(new_n439), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n249), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n470), .A2(new_n249), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n473), .B1(new_n571), .B2(new_n477), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT75), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n569), .A2(new_n485), .A3(new_n565), .A4(new_n566), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n574), .B2(new_n251), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(G200), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT6), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n579), .A2(new_n486), .A3(G107), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n582), .A2(new_n210), .B1(new_n206), .B2(new_n424), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n436), .B1(new_n401), .B2(new_n402), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n268), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n264), .A2(G97), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n504), .B2(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(G190), .B2(new_n575), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n574), .A2(new_n251), .ZN(new_n590));
  INV_X1    g0390(.A(new_n572), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n449), .B1(new_n585), .B2(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n575), .A2(new_n298), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n578), .A2(new_n589), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n316), .A2(new_n318), .A3(G244), .A4(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n323), .C2(new_n219), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n251), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n249), .A2(G274), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n467), .A2(new_n221), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n467), .B1(new_n249), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(G179), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n449), .B2(new_n604), .ZN(new_n606));
  INV_X1    g0406(.A(new_n426), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n264), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n316), .A2(new_n318), .A3(new_n210), .A4(G68), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT77), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n257), .A2(KEYINPUT77), .A3(new_n210), .A4(G68), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n210), .B1(new_n320), .B2(new_n611), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT76), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G97), .A2(G107), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n220), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n615), .B2(new_n618), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n613), .B(new_n614), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  AOI211_X1 g0421(.A(KEYINPUT78), .B(new_n608), .C1(new_n621), .C2(new_n268), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT78), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n609), .A2(new_n610), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n612), .A2(new_n611), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n614), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n619), .A2(new_n620), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n268), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n608), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n492), .A2(new_n426), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n606), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n492), .A2(new_n220), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n604), .B2(G200), .ZN(new_n635));
  OAI211_X1 g0435(.A(KEYINPUT79), .B(new_n635), .C1(new_n622), .C2(new_n630), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n602), .A2(new_n249), .ZN(new_n637));
  INV_X1    g0437(.A(new_n467), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n600), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n598), .B2(new_n251), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G190), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n624), .A2(new_n614), .A3(new_n625), .ZN(new_n643));
  INV_X1    g0443(.A(new_n620), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n615), .A2(new_n618), .A3(new_n616), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n304), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT78), .B1(new_n647), .B2(new_n608), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n628), .A2(new_n623), .A3(new_n629), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT79), .B1(new_n650), .B2(new_n635), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n595), .B(new_n633), .C1(new_n642), .C2(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n457), .A2(new_n564), .A3(new_n652), .ZN(G372));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n420), .B2(new_n421), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT18), .ZN(new_n656));
  INV_X1    g0456(.A(new_n356), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n367), .A2(new_n368), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n202), .B1(new_n402), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n406), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n304), .B1(new_n660), .B2(KEYINPUT16), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n661), .B2(new_n407), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n384), .A2(new_n389), .A3(G179), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n449), .B1(new_n384), .B2(new_n389), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n656), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n379), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(KEYINPUT88), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n454), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n314), .B1(new_n348), .B2(G190), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT71), .B1(new_n335), .B2(G200), .ZN(new_n671));
  INV_X1    g0471(.A(new_n350), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n343), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n655), .B(new_n668), .C1(new_n674), .C2(new_n411), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n295), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n301), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n575), .A2(G190), .ZN(new_n678));
  INV_X1    g0478(.A(new_n588), .ZN(new_n679));
  OAI21_X1  g0479(.A(G200), .B1(new_n575), .B2(new_n576), .ZN(new_n680));
  AOI211_X1 g0480(.A(KEYINPUT75), .B(new_n572), .C1(new_n574), .C2(new_n251), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n593), .A2(new_n594), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n550), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n634), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n622), .B2(new_n630), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT86), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(KEYINPUT86), .B(new_n685), .C1(new_n622), .C2(new_n630), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n604), .A2(G200), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n641), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n684), .A2(new_n633), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n561), .B1(new_n483), .B2(new_n556), .ZN(new_n694));
  AOI211_X1 g0494(.A(KEYINPUT21), .B(new_n555), .C1(new_n476), .C2(new_n482), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n553), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT87), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(KEYINPUT87), .B(new_n553), .C1(new_n694), .C2(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n523), .A2(new_n535), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n693), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n683), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n704), .B(new_n633), .C1(new_n642), .C2(new_n651), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT26), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n692), .A2(new_n707), .A3(new_n704), .A4(new_n633), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n633), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n677), .B1(new_n457), .B2(new_n710), .ZN(G369));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT89), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n716));
  INV_X1    g0516(.A(G213), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G343), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT90), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n495), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n698), .A2(new_n699), .A3(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n502), .B(new_n563), .C1(new_n495), .C2(new_n723), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n712), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n551), .B1(new_n523), .B2(new_n723), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n721), .B(KEYINPUT90), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n701), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n563), .A2(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n551), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n701), .A2(new_n723), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(G399));
  NAND3_X1  g0537(.A1(new_n213), .A2(KEYINPUT92), .A3(new_n245), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT92), .B1(new_n213), .B2(new_n245), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n618), .A2(G116), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT91), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(G1), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n217), .B2(new_n742), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n708), .A2(new_n633), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n701), .B1(new_n698), .B2(new_n699), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n749), .B(new_n706), .C1(new_n750), .C2(new_n693), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT29), .B1(new_n751), .B2(new_n723), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n536), .A2(new_n545), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n696), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n633), .B1(new_n754), .B2(new_n693), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n705), .A2(new_n707), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n692), .A2(KEYINPUT26), .A3(new_n704), .A4(new_n633), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n723), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT93), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n523), .A2(new_n503), .A3(new_n535), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT84), .B1(new_n537), .B2(new_n544), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n764), .B(new_n553), .C1(new_n694), .C2(new_n695), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n692), .A2(new_n633), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(new_n766), .A3(new_n684), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n756), .A2(new_n757), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n767), .A2(new_n768), .A3(new_n633), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT93), .A3(new_n723), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n752), .B1(new_n771), .B2(KEYINPUT29), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n652), .A2(new_n729), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n773), .A2(new_n551), .A3(new_n502), .A4(new_n563), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT30), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n465), .A2(new_n575), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n640), .A2(new_n531), .A3(new_n529), .A4(new_n552), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n552), .A2(new_n531), .A3(new_n529), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n604), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n780), .A2(KEYINPUT30), .A3(new_n465), .A4(new_n575), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(G179), .B1(new_n599), .B2(new_n603), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n592), .A2(new_n532), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n476), .B2(new_n482), .ZN(new_n785));
  OAI211_X1 g0585(.A(KEYINPUT31), .B(new_n729), .C1(new_n782), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n532), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n575), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n557), .B2(new_n558), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(new_n778), .A3(new_n781), .ZN(new_n791));
  AOI21_X1  g0591(.A(KEYINPUT31), .B1(new_n791), .B2(new_n729), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n712), .B1(new_n774), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n772), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n748), .B1(new_n795), .B2(G1), .ZN(G364));
  INV_X1    g0596(.A(G13), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n209), .B1(new_n798), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n741), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n727), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n725), .A2(new_n712), .A3(new_n726), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n725), .A2(new_n726), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n267), .B1(G20), .B2(new_n449), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT95), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n240), .A2(G45), .ZN(new_n812));
  INV_X1    g0612(.A(new_n213), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n257), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G45), .C2(new_n217), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n213), .A2(new_n257), .ZN(new_n816));
  INV_X1    g0616(.A(G355), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(G116), .B2(new_n213), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT94), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n811), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n801), .ZN(new_n821));
  INV_X1    g0621(.A(new_n809), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n210), .A2(new_n291), .A3(G179), .A4(G190), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G179), .A2(G200), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n210), .B1(new_n825), .B2(G190), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n824), .A2(new_n436), .B1(new_n486), .B2(new_n826), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n210), .A2(new_n298), .A3(new_n390), .A4(G200), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n257), .B1(new_n829), .B2(new_n201), .ZN(new_n830));
  NAND3_X1  g0630(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(G190), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n827), .B(new_n830), .C1(G68), .C2(new_n832), .ZN(new_n833));
  NOR4_X1   g0633(.A1(new_n210), .A2(new_n390), .A3(new_n291), .A4(G179), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n220), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n210), .A2(G190), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n825), .ZN(new_n838));
  INV_X1    g0638(.A(G159), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT32), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n831), .A2(new_n390), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n840), .A2(new_n841), .B1(new_n273), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n836), .B(new_n844), .C1(new_n841), .C2(new_n840), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n837), .A2(G179), .A3(new_n291), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n846), .A2(KEYINPUT96), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(KEYINPUT96), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n833), .B(new_n845), .C1(new_n206), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  INV_X1    g0651(.A(G329), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n846), .A2(new_n851), .B1(new_n838), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n257), .B(new_n853), .C1(G322), .C2(new_n828), .ZN(new_n854));
  INV_X1    g0654(.A(G317), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n855), .A2(KEYINPUT33), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(KEYINPUT33), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n832), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n826), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n834), .A2(G303), .B1(new_n859), .B2(G294), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n823), .A2(G283), .B1(G326), .B2(new_n842), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n854), .A2(new_n858), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n822), .B1(new_n850), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n820), .A2(new_n821), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n808), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n804), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G396));
  NAND2_X1  g0667(.A1(new_n729), .A2(new_n433), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n448), .A2(new_n454), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n454), .B2(new_n868), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n751), .B2(new_n723), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n723), .B(new_n870), .C1(new_n703), .C2(new_n709), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n794), .A3(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n642), .A2(new_n651), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n875), .A2(new_n595), .A3(new_n633), .A4(new_n723), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n793), .B1(new_n564), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(G330), .ZN(new_n878));
  INV_X1    g0678(.A(new_n873), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n874), .A2(new_n821), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n832), .ZN(new_n882));
  INV_X1    g0682(.A(G150), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(G143), .ZN(new_n885));
  INV_X1    g0685(.A(G137), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n829), .A2(new_n885), .B1(new_n886), .B2(new_n843), .ZN(new_n887));
  INV_X1    g0687(.A(new_n849), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n884), .B(new_n887), .C1(new_n888), .C2(G159), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n889), .A2(KEYINPUT34), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(KEYINPUT34), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n824), .A2(new_n202), .ZN(new_n892));
  INV_X1    g0692(.A(G132), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n257), .B1(new_n893), .B2(new_n838), .C1(new_n835), .C2(new_n273), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n892), .B(new_n894), .C1(G58), .C2(new_n859), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n890), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G283), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n835), .A2(new_n436), .B1(new_n897), .B2(new_n882), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(G303), .B2(new_n842), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n888), .A2(G116), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n367), .B1(new_n838), .B2(new_n851), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(G294), .B2(new_n828), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n859), .A2(G97), .B1(new_n823), .B2(G87), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n899), .A2(new_n900), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n822), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n809), .A2(new_n805), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n821), .B(new_n905), .C1(new_n206), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n870), .B2(new_n806), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n881), .A2(new_n908), .ZN(G384));
  INV_X1    g0709(.A(new_n582), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n493), .B(new_n216), .C1(new_n910), .C2(KEYINPUT35), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(KEYINPUT35), .B2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n358), .A2(new_n360), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n203), .A2(G50), .A3(G77), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(G50), .B2(new_n202), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G1), .A3(new_n797), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT97), .Z(new_n919));
  INV_X1    g0719(.A(new_n633), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n684), .A2(new_n633), .A3(new_n692), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n765), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n760), .B(new_n729), .C1(new_n922), .C2(new_n768), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT93), .B1(new_n769), .B2(new_n723), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT29), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n457), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT29), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n710), .B2(new_n729), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n929), .A2(new_n677), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n669), .A2(new_n723), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n873), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n402), .A2(new_n658), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G68), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT16), .B1(new_n934), .B2(new_n362), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n356), .B1(new_n371), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n936), .A2(new_n720), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n411), .B2(new_n422), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT100), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT37), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n379), .B2(new_n393), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n665), .A2(new_n719), .B1(new_n408), .B2(new_n356), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT99), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n417), .A2(new_n418), .A3(new_n719), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n379), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n408), .B(new_n356), .C1(new_n391), .C2(new_n392), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT99), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n940), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n936), .A2(new_n944), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n940), .B1(new_n950), .B2(new_n946), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n939), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  AOI211_X1 g0753(.A(KEYINPUT100), .B(new_n951), .C1(new_n943), .C2(new_n948), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n938), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT38), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(KEYINPUT38), .B(new_n938), .C1(new_n953), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n723), .A2(new_n345), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT14), .B1(new_n348), .B2(new_n449), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(new_n340), .A3(new_n339), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n351), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n729), .A2(new_n314), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n342), .A2(new_n673), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT98), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT98), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n960), .C1(new_n351), .C2(new_n962), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n932), .A2(new_n959), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT37), .B1(new_n662), .B2(new_n397), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n947), .B1(new_n972), .B2(new_n945), .ZN(new_n973));
  INV_X1    g0773(.A(new_n948), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n952), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT100), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n949), .A2(new_n939), .A3(new_n952), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT102), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT38), .A4(new_n938), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT39), .ZN(new_n981));
  INV_X1    g0781(.A(new_n958), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n719), .B1(new_n408), .B2(new_n356), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n655), .A2(new_n668), .A3(new_n410), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT101), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n946), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n654), .B1(new_n662), .B2(new_n665), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n662), .A2(KEYINPUT101), .A3(new_n397), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n379), .A2(KEYINPUT88), .A3(new_n419), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT37), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n983), .A2(new_n984), .B1(new_n991), .B2(new_n949), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT102), .B1(new_n992), .B2(KEYINPUT38), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n980), .B(new_n981), .C1(new_n982), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n343), .A2(new_n723), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n957), .A2(KEYINPUT39), .A3(new_n958), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n655), .A2(new_n668), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n719), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n971), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n930), .B(new_n1001), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n926), .A2(new_n877), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n966), .A2(new_n870), .A3(new_n968), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n1004), .A2(new_n877), .A3(KEYINPUT40), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n984), .A2(new_n983), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n990), .A2(KEYINPUT37), .B1(new_n943), .B2(new_n948), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n956), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n958), .A3(KEYINPUT102), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n1005), .A2(new_n1009), .A3(new_n980), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n966), .A2(new_n870), .A3(new_n968), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n774), .B2(new_n793), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT40), .B1(new_n959), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1003), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT38), .B1(new_n978), .B2(new_n938), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1012), .B1(new_n1015), .B2(new_n982), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT40), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1005), .A2(new_n1009), .A3(new_n980), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n926), .A3(new_n877), .A4(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1014), .A2(new_n1020), .A3(G330), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1002), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n209), .B2(new_n798), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1002), .A2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n919), .B1(new_n1023), .B2(new_n1024), .ZN(G367));
  OAI21_X1  g0825(.A(new_n595), .B1(new_n679), .B2(new_n723), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n704), .A2(new_n729), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n734), .A2(new_n735), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT105), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT105), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n734), .A2(new_n1031), .A3(new_n735), .A4(new_n1028), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT44), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n736), .B2(new_n1028), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n734), .A2(new_n735), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1038), .A2(KEYINPUT44), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1030), .A2(KEYINPUT45), .A3(new_n1032), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1035), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n732), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n734), .B1(new_n731), .B2(new_n733), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT106), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT107), .B1(new_n727), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1047), .B(new_n1049), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1035), .A2(new_n1040), .A3(new_n732), .A4(new_n1041), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n795), .A2(new_n1044), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1052), .A2(new_n795), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n741), .B(KEYINPUT41), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n799), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n733), .A2(new_n551), .A3(new_n1028), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(KEYINPUT42), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT104), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n753), .A2(new_n682), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n729), .B1(new_n1059), .B2(new_n683), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1056), .B2(KEYINPUT42), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n723), .B1(new_n688), .B2(new_n689), .ZN(new_n1063));
  MUX2_X1   g0863(.A(new_n766), .B(new_n920), .S(new_n1063), .Z(new_n1064));
  AND2_X1   g0864(.A1(new_n1064), .A2(KEYINPUT43), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1064), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT103), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1066), .A2(KEYINPUT103), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1068), .A2(KEYINPUT43), .A3(new_n1069), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n1062), .A2(new_n1065), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1072));
  AND4_X1   g0872(.A1(new_n1043), .A2(new_n1071), .A3(new_n1028), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1071), .A2(new_n1072), .B1(new_n1043), .B2(new_n1028), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1055), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n814), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n810), .B1(new_n213), .B2(new_n426), .C1(new_n1077), .C2(new_n235), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n801), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT108), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n838), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G137), .A2(new_n1081), .B1(new_n828), .B2(G150), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n201), .B2(new_n835), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n888), .B2(G50), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n826), .A2(new_n202), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n843), .A2(new_n885), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G159), .C2(new_n832), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n367), .B1(new_n823), .B2(G77), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT109), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n888), .A2(G283), .ZN(new_n1091));
  INV_X1    g0891(.A(G303), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n367), .B1(new_n829), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G317), .B2(new_n1081), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n824), .A2(new_n486), .B1(new_n851), .B2(new_n843), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n882), .A2(new_n527), .B1(new_n826), .B2(new_n436), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n834), .A2(G116), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT46), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1090), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT110), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT47), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n809), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n807), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1080), .B1(new_n1105), .B2(new_n1106), .C1(new_n1064), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1076), .A2(new_n1108), .ZN(G387));
  NAND3_X1  g0909(.A1(new_n728), .A2(new_n730), .A3(new_n807), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n814), .B1(new_n232), .B2(new_n246), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n745), .B2(new_n816), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n278), .A2(new_n273), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT50), .Z(new_n1114));
  AOI21_X1  g0914(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n745), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1112), .A2(new_n1116), .B1(new_n436), .B2(new_n813), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n801), .B1(new_n1117), .B2(new_n811), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n846), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1119), .A2(G68), .B1(new_n278), .B2(new_n832), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT111), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n257), .B1(new_n838), .B2(new_n883), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G50), .B2(new_n828), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n835), .A2(new_n206), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G97), .B2(new_n823), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n859), .A2(new_n607), .B1(G159), .B2(new_n842), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n257), .B1(new_n1081), .B2(G326), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n835), .A2(new_n527), .B1(new_n897), .B2(new_n826), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n828), .A2(G317), .B1(G311), .B2(new_n832), .ZN(new_n1130));
  INV_X1    g0930(.A(G322), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n843), .C1(new_n849), .C2(new_n1092), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT48), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1133), .B2(new_n1132), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT49), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1128), .B1(new_n493), .B2(new_n824), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1127), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1118), .B1(new_n1139), .B2(new_n809), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1050), .A2(new_n800), .B1(new_n1110), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n795), .A2(new_n1050), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n741), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n795), .A2(new_n1050), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(G393));
  NAND2_X1  g0945(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n741), .A3(new_n1052), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT113), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(KEYINPUT113), .A3(new_n741), .A4(new_n1052), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(KEYINPUT112), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT112), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1044), .A2(new_n1154), .A3(new_n1051), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n800), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n814), .A2(new_n243), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n807), .B(new_n809), .C1(new_n813), .C2(G97), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n821), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n849), .A2(new_n355), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n257), .B1(new_n885), .B2(new_n838), .C1(new_n824), .C2(new_n220), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n826), .A2(new_n206), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n835), .A2(new_n202), .B1(new_n273), .B2(new_n882), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n828), .A2(G159), .B1(G150), .B2(new_n842), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT51), .Z(new_n1166));
  AOI22_X1  g0966(.A1(new_n828), .A2(G311), .B1(G317), .B2(new_n842), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT52), .Z(new_n1168));
  OAI22_X1  g0968(.A1(new_n835), .A2(new_n897), .B1(new_n493), .B2(new_n826), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n367), .B1(new_n838), .B2(new_n1131), .C1(new_n527), .C2(new_n846), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n824), .A2(new_n436), .B1(new_n1092), .B2(new_n882), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1164), .A2(new_n1166), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1159), .B1(new_n822), .B2(new_n1173), .C1(new_n1028), .C2(new_n1107), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1156), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n1176), .ZN(G390));
  NAND3_X1  g0977(.A1(new_n794), .A2(new_n870), .A3(new_n970), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1009), .A2(new_n980), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n995), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n870), .B1(new_n923), .B2(new_n924), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n931), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n1183), .B2(new_n970), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n932), .A2(new_n970), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(new_n995), .B1(new_n997), .B2(new_n994), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n994), .A2(new_n997), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n969), .B1(new_n873), .B2(new_n931), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n996), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n969), .B1(new_n1182), .B2(new_n931), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1178), .C1(new_n1191), .C2(new_n1181), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1187), .A2(new_n800), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1188), .A2(new_n805), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n821), .B1(new_n355), .B2(new_n906), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n882), .A2(new_n886), .B1(new_n826), .B2(new_n839), .ZN(new_n1196));
  INV_X1    g0996(.A(G125), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n829), .A2(new_n893), .B1(new_n838), .B2(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G128), .C2(new_n842), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n367), .B1(new_n823), .B2(G50), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT116), .Z(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT53), .B1(new_n835), .B2(new_n883), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n883), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT54), .B(G143), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n888), .B2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1162), .B1(new_n832), .B2(G107), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n897), .B2(new_n843), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n367), .B1(new_n838), .B2(new_n527), .C1(new_n829), .C2(new_n493), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1210), .A2(new_n836), .A3(new_n892), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n486), .B2(new_n849), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1213), .A2(KEYINPUT117), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT117), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n809), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1194), .B(new_n1195), .C1(new_n1214), .C2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1193), .A2(KEYINPUT118), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT118), .B1(new_n1193), .B2(new_n1217), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n870), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n969), .B1(new_n878), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1178), .A2(new_n1223), .B1(new_n873), .B2(new_n931), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n931), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n771), .B2(new_n870), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1178), .A2(new_n1223), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1224), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n926), .A2(new_n794), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n929), .A2(new_n677), .A3(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1187), .A2(new_n1232), .A3(new_n1192), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1233), .A2(new_n741), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT114), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1227), .A2(new_n932), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1183), .B2(new_n1227), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT114), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n930), .A2(new_n1237), .A3(new_n1238), .A4(new_n1230), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n995), .B(new_n1180), .C1(new_n1226), .C2(new_n969), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1178), .B1(new_n1240), .B2(new_n1190), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1192), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1235), .B(new_n1239), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT115), .B1(new_n1234), .B2(new_n1243), .ZN(new_n1244));
  AND4_X1   g1044(.A1(KEYINPUT115), .A2(new_n1243), .A3(new_n741), .A4(new_n1233), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1221), .B1(new_n1244), .B2(new_n1245), .ZN(G378));
  NOR3_X1   g1046(.A1(new_n1010), .A2(new_n1013), .A3(new_n712), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1001), .A2(new_n1247), .A3(KEYINPUT121), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n287), .A2(new_n719), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n302), .B(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1250), .B(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1018), .A2(G330), .A3(new_n1019), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT121), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1018), .A2(KEYINPUT121), .A3(G330), .A4(new_n1019), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1256), .A2(new_n971), .A3(new_n998), .A4(new_n1000), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1248), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1255), .B1(new_n1248), .B2(new_n1257), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(new_n805), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n257), .A2(G41), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n897), .B2(new_n838), .C1(new_n829), .C2(new_n436), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n824), .A2(new_n201), .B1(new_n493), .B2(new_n843), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1085), .A4(new_n1124), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n882), .A2(new_n486), .B1(new_n846), .B2(new_n426), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT119), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT120), .Z(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(KEYINPUT58), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(KEYINPUT58), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G33), .A2(G41), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1262), .A2(G50), .A3(new_n1272), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n882), .A2(new_n893), .B1(new_n843), .B2(new_n1197), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G150), .B2(new_n859), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1119), .A2(G137), .B1(new_n828), .B2(G128), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(new_n835), .C2(new_n1204), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT59), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1081), .A2(G124), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1279), .B(new_n1272), .C1(new_n839), .C2(new_n824), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1277), .B2(KEYINPUT59), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1273), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1270), .A2(new_n1271), .A3(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1283), .A2(new_n809), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n821), .B(new_n1284), .C1(new_n273), .C2(new_n906), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1260), .A2(new_n800), .B1(new_n1261), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1231), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1233), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1248), .A2(new_n1257), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1255), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1248), .A2(new_n1257), .A3(new_n1255), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(KEYINPUT57), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n741), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1233), .A2(new_n1287), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1286), .B1(new_n1294), .B2(new_n1296), .ZN(G375));
  AOI21_X1  g1097(.A(new_n821), .B1(new_n202), .B2(new_n906), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n824), .A2(new_n206), .B1(new_n426), .B2(new_n826), .ZN(new_n1299));
  OAI221_X1 g1099(.A(new_n367), .B1(new_n838), .B2(new_n1092), .C1(new_n829), .C2(new_n897), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n1299), .B(new_n1300), .C1(new_n888), .C2(G107), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n835), .A2(new_n486), .B1(new_n527), .B2(new_n843), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(G116), .B2(new_n832), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n843), .A2(new_n893), .B1(new_n826), .B2(new_n273), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(G159), .B2(new_n834), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1119), .A2(G150), .B1(new_n1081), .B2(G128), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n367), .B1(new_n828), .B2(G137), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n832), .A2(new_n1205), .B1(new_n823), .B2(G58), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1301), .A2(new_n1303), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1310));
  OAI221_X1 g1110(.A(new_n1298), .B1(new_n822), .B2(new_n1310), .C1(new_n970), .C2(new_n806), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1229), .B2(new_n799), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT122), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT122), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1314), .B(new_n1311), .C1(new_n1229), .C2(new_n799), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1054), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1239), .A2(new_n1235), .A3(new_n1317), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(G381));
  OAI211_X1 g1120(.A(new_n866), .B(new_n1141), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(G387), .A2(G384), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1261), .A2(new_n1285), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1323), .B1(new_n1324), .B2(new_n799), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1260), .A2(new_n1295), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT57), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1258), .A2(new_n1259), .A3(new_n1327), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n742), .B1(new_n1329), .B2(new_n1295), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1325), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1243), .A2(new_n741), .A3(new_n1233), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1193), .A2(new_n1217), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT118), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1332), .A2(new_n1335), .A3(new_n1218), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(G390), .A2(G381), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1322), .A2(new_n1331), .A3(new_n1336), .A4(new_n1337), .ZN(G407));
  NOR2_X1   g1138(.A1(new_n717), .A2(G343), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(KEYINPUT123), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1331), .A2(new_n1336), .A3(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(G407), .A2(G213), .A3(new_n1341), .ZN(G409));
  AND3_X1   g1142(.A1(new_n1260), .A2(new_n1295), .A3(new_n1317), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1221), .B(new_n1332), .C1(new_n1343), .C2(new_n1325), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1335), .A2(new_n1218), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT115), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1332), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1234), .A2(KEYINPUT115), .A3(new_n1243), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1345), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1344), .B1(new_n1349), .B2(G375), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1339), .ZN(new_n1351));
  OAI21_X1  g1151(.A(KEYINPUT60), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1318), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT60), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1353), .B(new_n741), .C1(new_n1354), .C2(new_n1318), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1356), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1358), .A2(new_n1360), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1355), .A2(new_n1357), .A3(new_n1359), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1350), .A2(new_n1351), .A3(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1340), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1350), .A2(KEYINPUT62), .A3(new_n1363), .A4(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1366), .A2(new_n1368), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1355), .A2(new_n1357), .A3(new_n1359), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1359), .B1(new_n1355), .B2(new_n1357), .ZN(new_n1371));
  INV_X1    g1171(.A(G2897), .ZN(new_n1372));
  OAI22_X1  g1172(.A1(new_n1370), .A2(new_n1371), .B1(new_n1372), .B2(new_n1351), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1367), .A2(new_n1372), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1361), .A2(new_n1362), .A3(new_n1374), .ZN(new_n1375));
  AND2_X1   g1175(.A1(new_n1373), .A2(new_n1375), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1286), .B1(new_n1054), .B2(new_n1326), .ZN(new_n1377));
  AOI22_X1  g1177(.A1(G378), .A2(new_n1331), .B1(new_n1336), .B2(new_n1377), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1376), .B1(new_n1378), .B2(new_n1340), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT61), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1379), .A2(KEYINPUT127), .A3(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT127), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1373), .A2(new_n1375), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1383), .B1(new_n1350), .B2(new_n1367), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1382), .B1(new_n1384), .B2(KEYINPUT61), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1369), .A2(new_n1381), .A3(new_n1385), .ZN(new_n1386));
  AOI21_X1  g1186(.A(new_n1175), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(G393), .A2(G396), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1388), .A2(new_n1321), .ZN(new_n1389));
  AND2_X1   g1189(.A1(new_n1387), .A2(new_n1389), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1387), .A2(new_n1389), .ZN(new_n1391));
  OAI21_X1  g1191(.A(G387), .B1(new_n1390), .B2(new_n1391), .ZN(new_n1392));
  INV_X1    g1192(.A(new_n1389), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(G390), .A2(new_n1393), .ZN(new_n1394));
  AND2_X1   g1194(.A1(new_n1076), .A2(new_n1108), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1387), .A2(new_n1389), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1394), .A2(new_n1395), .A3(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1392), .A2(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1386), .A2(new_n1398), .ZN(new_n1399));
  INV_X1    g1199(.A(KEYINPUT126), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1376), .B1(new_n1378), .B2(new_n1339), .ZN(new_n1401));
  AND2_X1   g1201(.A1(new_n1363), .A2(KEYINPUT63), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1350), .A2(new_n1402), .A3(new_n1367), .ZN(new_n1403));
  AND3_X1   g1203(.A1(new_n1392), .A2(new_n1380), .A3(new_n1397), .ZN(new_n1404));
  NAND3_X1  g1204(.A1(new_n1401), .A2(new_n1403), .A3(new_n1404), .ZN(new_n1405));
  XNOR2_X1  g1205(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1406));
  INV_X1    g1206(.A(new_n1406), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(G378), .A2(new_n1331), .ZN(new_n1408));
  AOI21_X1  g1208(.A(new_n1339), .B1(new_n1408), .B2(new_n1344), .ZN(new_n1409));
  AOI21_X1  g1209(.A(new_n1407), .B1(new_n1409), .B2(new_n1363), .ZN(new_n1410));
  OAI21_X1  g1210(.A(new_n1400), .B1(new_n1405), .B2(new_n1410), .ZN(new_n1411));
  NAND3_X1  g1211(.A1(new_n1392), .A2(new_n1397), .A3(new_n1380), .ZN(new_n1412));
  NAND2_X1  g1212(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1413));
  AOI21_X1  g1213(.A(new_n1412), .B1(new_n1413), .B2(new_n1376), .ZN(new_n1414));
  NAND2_X1  g1214(.A1(new_n1364), .A2(new_n1406), .ZN(new_n1415));
  NAND4_X1  g1215(.A1(new_n1414), .A2(KEYINPUT126), .A3(new_n1415), .A4(new_n1403), .ZN(new_n1416));
  NAND2_X1  g1216(.A1(new_n1411), .A2(new_n1416), .ZN(new_n1417));
  NAND2_X1  g1217(.A1(new_n1399), .A2(new_n1417), .ZN(G405));
  NAND2_X1  g1218(.A1(G375), .A2(new_n1336), .ZN(new_n1419));
  AND2_X1   g1219(.A1(new_n1408), .A2(new_n1419), .ZN(new_n1420));
  XNOR2_X1  g1220(.A(new_n1420), .B(new_n1398), .ZN(new_n1421));
  INV_X1    g1221(.A(new_n1363), .ZN(new_n1422));
  XNOR2_X1  g1222(.A(new_n1421), .B(new_n1422), .ZN(G402));
endmodule


