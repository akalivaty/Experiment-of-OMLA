//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n452), .A2(G567), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT65), .Z(new_n456));
  AOI21_X1  g031(.A(new_n456), .B1(new_n451), .B2(G2106), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n465), .B2(G101), .ZN(new_n466));
  AND4_X1   g041(.A1(new_n463), .A2(new_n458), .A3(G101), .A4(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n464), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n469), .B1(new_n471), .B2(new_n459), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT66), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G113), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g055(.A(KEYINPUT67), .B(G2105), .C1(new_n472), .C2(new_n477), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n468), .B1(new_n480), .B2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n471), .A2(new_n459), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n458), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n471), .B2(new_n459), .ZN(new_n495));
  AND2_X1   g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n458), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n471), .B2(new_n459), .ZN(new_n499));
  AND2_X1   g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  OAI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(KEYINPUT71), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n514), .B2(KEYINPUT71), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI211_X1 g096(.A(G50), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(KEYINPUT69), .A3(G50), .A4(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n516), .A2(G88), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n507), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n520), .A2(new_n521), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n534), .B2(new_n511), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G88), .B1(new_n524), .B2(new_n526), .ZN(new_n536));
  INV_X1    g111(.A(G62), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n534), .B2(new_n511), .ZN(new_n538));
  INV_X1    g113(.A(new_n518), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n536), .A2(new_n540), .A3(KEYINPUT72), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(new_n541), .ZN(G166));
  NAND2_X1  g117(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n534), .A2(new_n544), .A3(new_n511), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n546), .A2(G63), .A3(G651), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n531), .A2(new_n510), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G51), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n516), .A2(new_n525), .ZN(new_n552));
  INV_X1    g127(.A(G89), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n549), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n547), .A2(new_n554), .ZN(G168));
  AOI22_X1  g130(.A1(new_n546), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n508), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n535), .A2(G90), .B1(new_n548), .B2(G52), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  AOI22_X1  g135(.A1(new_n546), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n508), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT74), .B(G43), .Z(new_n563));
  AOI22_X1  g138(.A1(new_n535), .A2(G81), .B1(new_n548), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND3_X1  g147(.A1(new_n548), .A2(KEYINPUT76), .A3(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n552), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n508), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G299));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n536), .A2(new_n540), .A3(KEYINPUT72), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT72), .B1(new_n536), .B2(new_n540), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n530), .A2(new_n541), .A3(KEYINPUT77), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G303));
  AOI22_X1  g162(.A1(new_n535), .A2(G87), .B1(new_n548), .B2(G49), .ZN(new_n588));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n543), .A2(new_n589), .A3(new_n545), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n590), .A2(new_n591), .A3(G651), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n590), .B2(G651), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(new_n548), .A2(G48), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n552), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n516), .B2(G61), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT79), .B1(new_n601), .B2(G651), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n604));
  NOR3_X1   g179(.A1(new_n600), .A2(new_n604), .A3(new_n508), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n597), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G305));
  AOI22_X1  g183(.A1(new_n535), .A2(G85), .B1(new_n548), .B2(G47), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n546), .A2(G60), .ZN(new_n610));
  NAND2_X1  g185(.A1(G72), .A2(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT80), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n612), .A2(KEYINPUT80), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(new_n535), .A2(G92), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT10), .Z(new_n622));
  AOI22_X1  g197(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(new_n508), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G54), .B2(new_n548), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G171), .B2(new_n627), .ZN(G284));
  OAI21_X1  g204(.A(new_n628), .B1(G171), .B2(new_n627), .ZN(G321));
  NAND2_X1  g205(.A1(G286), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n579), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(new_n579), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G860), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n626), .B1(G559), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g211(.A1(new_n565), .A2(new_n627), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n626), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n483), .A2(new_n465), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT83), .B(G2100), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n485), .A2(G123), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n488), .A2(G135), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n458), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n645), .A2(new_n646), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2451), .B(G2454), .Z(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n667), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  INV_X1    g252(.A(new_n675), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(KEYINPUT85), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(KEYINPUT85), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n672), .B(KEYINPUT17), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n681), .C1(new_n678), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n674), .A3(new_n678), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(new_n652), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT86), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n693), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  AOI211_X1 g272(.A(new_n695), .B(new_n697), .C1(new_n690), .C2(new_n694), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1981), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n700), .B(new_n704), .ZN(G229));
  INV_X1    g280(.A(G290), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G16), .B2(G24), .ZN(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT88), .B(G29), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n485), .A2(G119), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n488), .A2(G131), .ZN(new_n716));
  OR2_X1    g291(.A1(G95), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n713), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NOR3_X1   g298(.A1(new_n710), .A2(new_n711), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G6), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n607), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT89), .Z(new_n730));
  MUX2_X1   g305(.A(G23), .B(G288), .S(G16), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT90), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT33), .B(G1976), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G22), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G166), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1971), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n730), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT34), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n724), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n725), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n566), .B2(new_n725), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G1341), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n712), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n485), .A2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n488), .A2(G140), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n458), .A2(G116), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n753), .A2(KEYINPUT91), .A3(G29), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT91), .B1(new_n753), .B2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n748), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n725), .A2(G4), .ZN(new_n759));
  INV_X1    g334(.A(new_n626), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n725), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n746), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n725), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  INV_X1    g345(.A(G32), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n488), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n485), .A2(G129), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(new_n771), .B(new_n777), .S(G29), .Z(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n713), .A2(G35), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n713), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT29), .B(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G11), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT30), .B(G28), .Z(new_n788));
  OAI221_X1 g363(.A(new_n787), .B1(G29), .B2(new_n788), .C1(new_n651), .C2(new_n712), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n780), .A2(new_n781), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n725), .A2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G168), .B2(new_n725), .ZN(new_n792));
  INV_X1    g367(.A(G1966), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n770), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G139), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n487), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n458), .B2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G33), .B(new_n803), .S(G29), .Z(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G2072), .ZN(new_n805));
  INV_X1    g380(.A(G2084), .ZN(new_n806));
  NAND2_X1  g381(.A1(G160), .A2(G29), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT24), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(G34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(G34), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n712), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n804), .A2(G2072), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n806), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT94), .Z(new_n815));
  NOR2_X1   g390(.A1(new_n713), .A2(G27), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G164), .B2(new_n713), .ZN(new_n817));
  INV_X1    g392(.A(G2078), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n805), .A2(new_n813), .A3(new_n815), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n725), .A2(G5), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G171), .B2(new_n725), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1961), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n795), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n743), .A2(new_n765), .A3(new_n766), .A4(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  NAND2_X1  g401(.A1(new_n760), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n546), .A2(G67), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n508), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n548), .A2(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n552), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n566), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n565), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n828), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n634), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n835), .A2(new_n634), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n753), .B(new_n505), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n803), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n776), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n485), .A2(G130), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n458), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G142), .B2(new_n488), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(new_n642), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n719), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n850), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(G160), .B(new_n651), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n492), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n860), .A2(KEYINPUT96), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT96), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  INV_X1    g441(.A(new_n862), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n858), .B(new_n867), .C1(KEYINPUT97), .C2(new_n859), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n859), .A2(KEYINPUT97), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g447(.A1(new_n837), .A2(new_n627), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n839), .B(new_n638), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n760), .B(new_n579), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n875), .B(KEYINPUT41), .Z(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(G288), .B(G166), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n706), .A2(KEYINPUT98), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n884));
  NAND2_X1  g459(.A1(G290), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(G305), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(G305), .B1(new_n883), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n881), .A3(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT99), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n880), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n873), .B1(new_n893), .B2(new_n627), .ZN(G295));
  OAI21_X1  g469(.A(new_n873), .B1(new_n893), .B2(new_n627), .ZN(G331));
  NAND2_X1  g470(.A1(G301), .A2(G168), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT100), .Z(new_n897));
  NOR2_X1   g472(.A1(G301), .A2(G168), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT101), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n839), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n839), .A3(new_n899), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n876), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n900), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n905), .B2(new_n878), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n889), .A2(new_n891), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n866), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n889), .B2(new_n891), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n889), .A2(new_n891), .ZN(new_n911));
  INV_X1    g486(.A(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n866), .A4(new_n907), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT44), .Z(G397));
  INV_X1    g492(.A(KEYINPUT126), .ZN(new_n918));
  NAND2_X1  g493(.A1(G160), .A2(G40), .ZN(new_n919));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n505), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(G290), .A2(G1986), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n776), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n753), .B(new_n757), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n719), .B(new_n722), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(KEYINPUT102), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(KEYINPUT102), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G290), .A2(G1986), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n925), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n505), .A2(new_n939), .A3(new_n920), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n505), .B2(new_n920), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT50), .ZN(new_n942));
  INV_X1    g517(.A(G40), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n943), .B(new_n468), .C1(new_n480), .C2(new_n481), .ZN(new_n944));
  INV_X1    g519(.A(new_n921), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2090), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n920), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n923), .A2(new_n944), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n737), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n938), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n938), .B1(KEYINPUT104), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n585), .A2(new_n586), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(KEYINPUT104), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n960));
  INV_X1    g535(.A(new_n958), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n585), .A2(new_n586), .A3(new_n961), .A4(new_n956), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n960), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n954), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1976), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT52), .B1(G288), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n940), .A2(new_n941), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n938), .B1(new_n968), .B2(new_n944), .ZN(new_n969));
  OAI211_X1 g544(.A(G1976), .B(new_n588), .C1(new_n592), .C2(new_n593), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n921), .A2(KEYINPUT103), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n505), .A2(new_n939), .A3(new_n920), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n944), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n974), .A3(G8), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT52), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1981), .ZN(new_n978));
  INV_X1    g553(.A(new_n597), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n979), .C1(new_n602), .C2(new_n605), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n600), .A2(new_n508), .ZN(new_n981));
  OAI21_X1  g556(.A(G1981), .B1(new_n981), .B2(new_n597), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT106), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(G1981), .C1(new_n981), .C2(new_n597), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n980), .A2(new_n983), .A3(KEYINPUT49), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n969), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(KEYINPUT107), .A3(new_n990), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n977), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n965), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n946), .B1(new_n972), .B2(new_n973), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(new_n919), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT109), .B(new_n944), .C1(new_n968), .C2(new_n946), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n945), .A2(new_n946), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n953), .B1(new_n1001), .B2(G2090), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n1002), .A2(G8), .B1(new_n959), .B2(new_n962), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT121), .B1(new_n995), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1961), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n942), .B2(new_n947), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n922), .B1(new_n940), .B2(new_n941), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n951), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n505), .A2(KEYINPUT110), .A3(KEYINPUT45), .A4(new_n920), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(G2078), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1007), .A2(new_n1011), .A3(new_n944), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n952), .B2(G2078), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1006), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G171), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(KEYINPUT118), .A3(G171), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1007), .A2(new_n1011), .A3(new_n944), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n793), .ZN(new_n1023));
  INV_X1    g598(.A(new_n942), .ZN(new_n1024));
  INV_X1    g599(.A(new_n947), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n806), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1026), .A3(G168), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n938), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT51), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1028), .B(KEYINPUT51), .C1(new_n1031), .C2(new_n1030), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT62), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(G286), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1002), .A2(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n959), .A2(new_n962), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n965), .A4(new_n994), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1004), .A2(new_n1021), .A3(new_n1037), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1030), .A2(G168), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1040), .A2(new_n1054), .A3(new_n965), .A4(new_n994), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n954), .B1(new_n959), .B2(new_n962), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n1056), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(new_n965), .A3(new_n994), .A4(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n991), .A2(new_n988), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n986), .A2(new_n969), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n993), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(new_n971), .A3(new_n976), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n965), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n969), .ZN(new_n1066));
  OR2_X1    g641(.A1(G288), .A2(G1976), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1069), .B2(new_n980), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT108), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n992), .B2(new_n993), .ZN(new_n1072));
  INV_X1    g647(.A(new_n980), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n969), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1039), .A2(KEYINPUT105), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n994), .A2(new_n1077), .A3(new_n954), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1057), .A2(new_n1060), .B1(new_n1071), .B2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1016), .A2(KEYINPUT118), .A3(G171), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT118), .B1(new_n1016), .B2(G171), .ZN(new_n1083));
  INV_X1    g658(.A(new_n468), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(G40), .A3(new_n478), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT119), .B1(new_n923), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT45), .B1(new_n505), .B2(new_n920), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1085), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n951), .B(new_n1013), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1091));
  AND4_X1   g666(.A1(G301), .A2(new_n1091), .A3(new_n1015), .A4(new_n1006), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1082), .A2(new_n1083), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n1093), .B2(KEYINPUT54), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1095), .B(new_n1096), .C1(new_n1021), .C2(new_n1092), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1006), .A2(new_n1015), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1099), .B2(new_n1091), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n1016), .B2(G171), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1029), .A2(new_n1032), .B1(G286), .B2(new_n1030), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1034), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1098), .A2(new_n1004), .A3(new_n1042), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1956), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1001), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n952), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT56), .B(G2072), .Z(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT112), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT111), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1113), .A2(KEYINPUT111), .ZN(new_n1115));
  NAND3_X1  g690(.A1(G299), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n579), .A2(KEYINPUT111), .A3(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT61), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n762), .B1(new_n942), .B2(new_n947), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n974), .A2(G2067), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n760), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1125), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n626), .B1(new_n1127), .B2(new_n1123), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT60), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n626), .A2(KEYINPUT60), .ZN(new_n1131));
  INV_X1    g706(.A(new_n974), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(G1341), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1132), .A2(new_n1134), .B1(G1996), .B2(new_n952), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n566), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(KEYINPUT59), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1130), .A2(new_n1131), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1137), .B2(KEYINPUT59), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n566), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1129), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1122), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1120), .A2(new_n1146), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1145), .A2(KEYINPUT61), .A3(new_n1119), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1128), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1119), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1144), .A2(new_n1148), .B1(new_n1121), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1081), .B1(new_n1105), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1045), .A2(new_n1053), .B1(new_n1152), .B2(KEYINPUT122), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1081), .B(new_n1154), .C1(new_n1105), .C2(new_n1151), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n937), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT48), .ZN(new_n1157));
  INV_X1    g732(.A(new_n926), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n925), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n926), .A2(KEYINPUT48), .A3(new_n924), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n924), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT46), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n925), .B2(G1996), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n924), .A2(KEYINPUT46), .A3(new_n927), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n929), .A2(new_n777), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1164), .B(new_n1165), .C1(new_n925), .C2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT125), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT47), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n720), .A2(new_n722), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n930), .A2(new_n1170), .B1(G2067), .B2(new_n753), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n924), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1162), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n918), .B1(new_n1156), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n1177), .A3(new_n1045), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1155), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n937), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1173), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT126), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1174), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g758(.A(G319), .B1(new_n669), .B2(new_n670), .ZN(new_n1185));
  NOR3_X1   g759(.A1(G229), .A2(G227), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g760(.A(new_n1186), .B1(new_n865), .B2(new_n870), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n910), .B2(new_n915), .ZN(new_n1188));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1189));
  XNOR2_X1  g763(.A(new_n1188), .B(new_n1189), .ZN(G308));
  XNOR2_X1  g764(.A(new_n1188), .B(KEYINPUT127), .ZN(G225));
endmodule


