//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G104), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n193), .A2(KEYINPUT77), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n195), .A2(new_n190), .A3(new_n194), .A4(new_n192), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n189), .A2(G104), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n194), .B1(new_n201), .B2(new_n192), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(KEYINPUT2), .B2(G113), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n206));
  INV_X1    g020(.A(G113), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT70), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT2), .A2(G113), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(KEYINPUT71), .A2(KEYINPUT2), .A3(G113), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n205), .A2(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G116), .B(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT5), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(KEYINPUT5), .A3(G119), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(new_n207), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n200), .A2(new_n203), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n195), .A2(new_n190), .A3(new_n192), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n199), .B2(new_n196), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n205), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n211), .A2(new_n212), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n214), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n213), .A2(new_n214), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n221), .A2(new_n232), .A3(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n220), .B1(new_n224), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n187), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n220), .B(new_n236), .C1(new_n224), .C2(new_n234), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT82), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n221), .A2(new_n232), .A3(G101), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n229), .B2(new_n230), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n232), .B1(new_n221), .B2(G101), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n197), .A2(new_n198), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n197), .A2(new_n198), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n202), .B1(new_n196), .B2(new_n199), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n243), .A2(new_n247), .B1(new_n248), .B2(new_n219), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n241), .B1(new_n249), .B2(new_n236), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n238), .B1(new_n240), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT83), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  XNOR2_X1  g068(.A(G143), .B(G146), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n257), .C2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G128), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT68), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT69), .B(new_n256), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(G146), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n255), .A2(KEYINPUT67), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT1), .B1(new_n257), .B2(G146), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(G128), .A3(new_n258), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT69), .B1(new_n276), .B2(new_n256), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n254), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n255), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT0), .B(G128), .Z(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n255), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G125), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT85), .B(G224), .Z(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(G953), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT84), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n284), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n235), .A2(new_n187), .A3(new_n237), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT83), .B(new_n238), .C1(new_n240), .C2(new_n250), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n253), .A2(new_n288), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n236), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n248), .A2(new_n219), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n220), .ZN(new_n296));
  INV_X1    g110(.A(new_n240), .ZN(new_n297));
  INV_X1    g111(.A(new_n250), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n284), .B(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G210), .B1(G237), .B2(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT87), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n291), .A2(new_n302), .A3(new_n305), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT91), .B1(new_n264), .B2(G143), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n257), .A3(G128), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n257), .A2(G128), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n216), .A2(G122), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n216), .A2(G122), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n189), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n321), .A3(G107), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT13), .B1(new_n312), .B2(new_n314), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(new_n317), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT92), .B1(new_n328), .B2(new_n316), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT13), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n315), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT13), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n318), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G134), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n325), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n315), .A2(new_n318), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G134), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n319), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n189), .B1(new_n320), .B2(KEYINPUT14), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(new_n322), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n322), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT9), .B(G234), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n345), .A2(new_n346), .A3(G953), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n336), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n325), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n333), .A2(new_n334), .A3(G134), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n334), .B1(new_n333), .B2(G134), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n347), .B1(new_n353), .B2(new_n343), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n311), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT93), .ZN(new_n356));
  INV_X1    g170(.A(G478), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT15), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n348), .B1(new_n336), .B2(new_n344), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n343), .A3(new_n347), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n311), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n358), .B(KEYINPUT94), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n311), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(G952), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(G902), .A3(G953), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT21), .B(G898), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n377));
  NOR2_X1   g191(.A1(G237), .A2(G953), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(G143), .A3(G214), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n378), .B2(G214), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT18), .B(G131), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G125), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n254), .A2(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n260), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n381), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n379), .A3(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n382), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT74), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT74), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n384), .A2(new_n385), .A3(new_n397), .A4(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n260), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT19), .B1(new_n384), .B2(new_n385), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT19), .ZN(new_n402));
  AOI21_X1  g216(.A(G146), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G131), .B1(new_n380), .B2(new_n381), .ZN(new_n405));
  INV_X1    g219(.A(G131), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n390), .A2(new_n406), .A3(new_n379), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n393), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n191), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT88), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT74), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n398), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G146), .ZN(new_n416));
  INV_X1    g230(.A(new_n402), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n260), .B1(new_n417), .B2(new_n400), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n408), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n382), .A2(new_n389), .A3(new_n392), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n405), .A2(new_n407), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n260), .B(new_n398), .C1(new_n413), .C2(new_n414), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n416), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT17), .B(G131), .C1(new_n380), .C2(new_n381), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n393), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n412), .A2(new_n423), .B1(new_n432), .B2(new_n411), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n377), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n429), .B(KEYINPUT89), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n411), .B(new_n420), .C1(new_n437), .C2(new_n427), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n421), .A2(new_n422), .ZN(new_n439));
  AOI211_X1 g253(.A(KEYINPUT88), .B(new_n411), .C1(new_n419), .C2(new_n420), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT90), .A3(new_n434), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n442), .A3(KEYINPUT20), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT90), .B1(new_n441), .B2(new_n434), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n420), .B1(new_n437), .B2(new_n427), .ZN(new_n446));
  INV_X1    g260(.A(new_n411), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n438), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n311), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n444), .A2(new_n445), .B1(G475), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n367), .A2(new_n376), .A3(new_n443), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n310), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G137), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n369), .A2(G221), .A3(G234), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n454), .B(new_n455), .Z(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n264), .A2(G119), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT24), .B(G110), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n458), .B2(G128), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n264), .A2(KEYINPUT23), .A3(G119), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n459), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(G110), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n426), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n399), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n461), .A2(new_n462), .ZN(new_n471));
  INV_X1    g285(.A(G110), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n465), .A2(new_n466), .A3(new_n472), .A4(new_n459), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n388), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n399), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n416), .A2(new_n388), .A3(new_n474), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT75), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n457), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n478), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(KEYINPUT75), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n470), .A4(new_n456), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n311), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT76), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n346), .B1(G234), .B2(new_n311), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n488), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT25), .A4(new_n311), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT76), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n482), .A2(new_n485), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n490), .A2(G902), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n491), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n378), .A2(G210), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT27), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT11), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n316), .B2(G137), .ZN(new_n506));
  INV_X1    g320(.A(G137), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT11), .A3(G134), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n316), .A2(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n510), .A2(KEYINPUT65), .A3(G131), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT65), .B1(new_n510), .B2(G131), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n506), .A2(new_n508), .A3(new_n406), .A4(new_n509), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n282), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n508), .A2(new_n509), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(new_n515), .A3(new_n406), .A4(new_n506), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(KEYINPUT64), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n521));
  XNOR2_X1  g335(.A(G134), .B(G137), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n406), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n316), .A2(G137), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n507), .A2(G134), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT66), .B(G131), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n519), .A2(new_n520), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n272), .B2(new_n277), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n231), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT72), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n225), .A2(new_n226), .A3(new_n214), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n214), .B1(new_n225), .B2(new_n226), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n517), .A3(new_n528), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n504), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n504), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n503), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n231), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n523), .A2(new_n526), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n514), .A2(KEYINPUT64), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n514), .A2(KEYINPUT64), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n277), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n263), .A2(new_n271), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n510), .A2(G131), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT65), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n510), .A2(KEYINPUT65), .A3(G131), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n519), .A2(new_n520), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n281), .A2(new_n255), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n280), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT30), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n517), .A2(new_n528), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n542), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n537), .A2(new_n502), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT31), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n517), .A2(new_n528), .A3(new_n559), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n559), .B1(new_n517), .B2(new_n528), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n231), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n537), .A4(new_n502), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n541), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(G472), .A2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT32), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT29), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n539), .A2(new_n502), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n538), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n502), .B1(new_n566), .B2(new_n537), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n531), .A2(new_n535), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n549), .A2(new_n557), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n542), .B1(new_n517), .B2(new_n528), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT28), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n503), .B1(new_n537), .B2(new_n504), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT29), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n503), .B1(new_n561), .B2(new_n583), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT73), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n578), .A2(new_n577), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n529), .A2(new_n582), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n537), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT28), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n581), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n498), .B1(new_n575), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G221), .B1(new_n345), .B2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n600));
  XNOR2_X1  g414(.A(G110), .B(G140), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n369), .A2(G227), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT80), .B1(new_n513), .B2(new_n516), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT78), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT67), .B1(new_n255), .B2(new_n265), .ZN(new_n607));
  AND4_X1   g421(.A1(KEYINPUT67), .A2(new_n265), .A3(new_n261), .A4(new_n266), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT78), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n273), .A2(G128), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n256), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n248), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n203), .B1(new_n245), .B2(new_n246), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n548), .A3(new_n547), .ZN(new_n616));
  AOI211_X1 g430(.A(KEYINPUT12), .B(new_n605), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT12), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n614), .ZN(new_n619));
  INV_X1    g433(.A(new_n605), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n282), .A2(new_n233), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n200), .B2(new_n244), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n614), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n554), .A2(KEYINPUT79), .A3(new_n555), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT79), .B1(new_n554), .B2(new_n555), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n248), .B(KEYINPUT10), .C1(new_n277), .C2(new_n272), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n604), .B1(new_n622), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n513), .A2(new_n516), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n626), .B2(new_n630), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n633), .A2(new_n635), .A3(new_n603), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n600), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n271), .A2(new_n606), .B1(new_n256), .B2(new_n611), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n615), .B1(new_n610), .B2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n248), .A2(new_n272), .A3(new_n277), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n620), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT12), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n619), .A2(new_n618), .A3(new_n620), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n603), .B1(new_n644), .B2(new_n633), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n626), .A2(new_n630), .ZN(new_n646));
  INV_X1    g460(.A(new_n634), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n631), .A3(new_n604), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(KEYINPUT81), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n637), .A2(G469), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G469), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n311), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n603), .B1(new_n633), .B2(new_n635), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n642), .A2(new_n631), .A3(new_n604), .A4(new_n643), .ZN(new_n655));
  AOI21_X1  g469(.A(G902), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n653), .B1(new_n656), .B2(new_n652), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n599), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n453), .A2(new_n597), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G101), .ZN(G3));
  NAND2_X1  g474(.A1(new_n569), .A2(new_n311), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n661), .A2(G472), .B1(new_n570), .B2(new_n569), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n658), .A2(new_n497), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n362), .B1(new_n361), .B2(new_n311), .ZN(new_n664));
  AOI211_X1 g478(.A(KEYINPUT93), .B(G902), .C1(new_n359), .C2(new_n360), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT95), .B1(new_n666), .B2(new_n357), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n356), .A2(KEYINPUT95), .A3(new_n357), .A4(new_n363), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n361), .A2(KEYINPUT33), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n361), .A2(KEYINPUT33), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n311), .A2(G478), .ZN(new_n673));
  OAI22_X1  g487(.A1(new_n667), .A2(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n451), .A2(new_n443), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n376), .A3(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n663), .A2(new_n310), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT34), .B(G104), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G6));
  AND3_X1   g493(.A1(new_n291), .A2(new_n302), .A3(new_n305), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n305), .B1(new_n291), .B2(new_n302), .ZN(new_n681));
  INV_X1    g495(.A(new_n308), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT97), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n364), .A2(new_n366), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n443), .A3(new_n451), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n375), .B(KEYINPUT96), .Z(new_n688));
  NAND4_X1  g502(.A1(new_n683), .A2(new_n684), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n688), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT97), .B1(new_n690), .B2(new_n686), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n663), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT35), .B(G107), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  NAND2_X1  g508(.A1(new_n491), .A2(new_n494), .ZN(new_n695));
  OR4_X1    g509(.A1(KEYINPUT36), .A2(new_n479), .A3(new_n481), .A4(new_n457), .ZN(new_n696));
  OAI22_X1  g510(.A1(new_n479), .A2(new_n481), .B1(KEYINPUT36), .B2(new_n457), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n696), .A2(new_n496), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n453), .A2(new_n658), .A3(new_n662), .A4(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  AND2_X1   g517(.A1(new_n451), .A2(new_n443), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT98), .ZN(new_n705));
  INV_X1    g519(.A(G900), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n371), .B1(new_n373), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n704), .A2(new_n705), .A3(new_n685), .A4(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n685), .A2(new_n443), .A3(new_n451), .A4(new_n708), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT98), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n658), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n572), .A2(new_n574), .B1(new_n595), .B2(G472), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n698), .B1(new_n491), .B2(new_n494), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n310), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  NOR2_X1   g531(.A1(new_n680), .A2(new_n681), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n451), .A2(new_n443), .B1(new_n364), .B2(new_n366), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n720), .A2(new_n682), .A3(new_n700), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT100), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n561), .A2(new_n583), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n503), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n311), .B1(new_n592), .B2(new_n502), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n724), .B1(new_n575), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n573), .B1(new_n569), .B2(new_n570), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n728), .B(new_n724), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n707), .B(KEYINPUT39), .Z(new_n735));
  AOI21_X1  g549(.A(KEYINPUT40), .B1(new_n658), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n658), .A2(KEYINPUT40), .A3(new_n735), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n723), .B(new_n734), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G143), .ZN(G45));
  AOI21_X1  g553(.A(new_n714), .B1(new_n575), .B2(new_n596), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n673), .B1(new_n670), .B2(new_n671), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n356), .A2(new_n357), .A3(new_n363), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n744), .B2(new_n668), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n704), .A3(new_n707), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n683), .A3(new_n658), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  NOR3_X1   g562(.A1(new_n745), .A2(new_n704), .A3(new_n375), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n656), .A2(new_n652), .ZN(new_n750));
  INV_X1    g564(.A(new_n655), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n604), .B1(new_n648), .B2(new_n631), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n652), .B(new_n311), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n598), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n597), .A2(new_n683), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  AND3_X1   g572(.A1(new_n581), .A2(new_n589), .A3(new_n594), .ZN(new_n759));
  INV_X1    g573(.A(G472), .ZN(new_n760));
  OAI22_X1  g574(.A1(new_n759), .A2(new_n760), .B1(new_n730), .B2(new_n731), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n755), .A2(new_n761), .A3(new_n497), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n689), .B2(new_n691), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n216), .ZN(G18));
  NOR2_X1   g578(.A1(new_n754), .A2(new_n452), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n740), .A2(new_n765), .A3(new_n683), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT101), .B(G119), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G21));
  NAND2_X1  g582(.A1(new_n661), .A2(G472), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n563), .A2(new_n568), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n502), .B1(new_n593), .B2(new_n539), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n570), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n497), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n750), .A2(new_n598), .A3(new_n753), .A4(new_n688), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n307), .A2(new_n721), .A3(new_n308), .A4(new_n309), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NOR2_X1   g593(.A1(new_n310), .A2(new_n754), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n700), .A2(new_n769), .A3(new_n772), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n782), .A3(new_n746), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G125), .ZN(G27));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n682), .B1(new_n307), .B2(new_n309), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n645), .A2(G469), .A3(new_n649), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n599), .B1(new_n657), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n761), .A2(new_n786), .A3(new_n497), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n674), .A2(new_n675), .A3(new_n708), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n308), .B1(new_n680), .B2(new_n681), .ZN(new_n792));
  INV_X1    g606(.A(new_n653), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n753), .A2(new_n793), .A3(new_n787), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n598), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n597), .A3(KEYINPUT42), .A4(new_n746), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n791), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G131), .ZN(G33));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n597), .A3(new_n709), .A4(new_n711), .ZN(new_n800));
  XNOR2_X1  g614(.A(KEYINPUT102), .B(G134), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(G36));
  INV_X1    g616(.A(new_n753), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n637), .B2(new_n650), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n645), .A2(KEYINPUT45), .A3(new_n649), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(G469), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n793), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT46), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n598), .A3(new_n735), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n662), .A2(new_n714), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n675), .B(KEYINPUT103), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n674), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT43), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n745), .A2(KEYINPUT43), .A3(new_n675), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT104), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n815), .A2(KEYINPUT104), .A3(new_n816), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n812), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n786), .B(new_n811), .C1(new_n821), .C2(KEYINPUT44), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(KEYINPUT44), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT105), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT105), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n825), .A3(KEYINPUT44), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n507), .ZN(G39));
  NOR4_X1   g642(.A1(new_n790), .A2(new_n761), .A3(new_n792), .A4(new_n497), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n810), .A2(new_n598), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(KEYINPUT47), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(KEYINPUT47), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT106), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT107), .B(G140), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(G42));
  NAND3_X1  g654(.A1(new_n497), .A2(new_n308), .A3(new_n598), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT108), .Z(new_n842));
  INV_X1    g656(.A(new_n814), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n656), .A2(new_n652), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n803), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT109), .Z(new_n848));
  INV_X1    g662(.A(new_n734), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n844), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n849), .A3(new_n720), .A4(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n675), .A2(new_n685), .A3(new_n707), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n740), .A2(new_n658), .A3(new_n786), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n796), .A2(new_n746), .A3(new_n782), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n800), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(new_n798), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT110), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n761), .A2(new_n658), .A3(new_n497), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n675), .A2(new_n685), .A3(new_n375), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n683), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n718), .A2(new_n859), .A3(new_n308), .A4(new_n700), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n651), .A2(new_n657), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n662), .A3(new_n598), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n858), .A2(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n686), .B1(new_n745), .B2(new_n704), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n683), .A3(new_n688), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n663), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n857), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n863), .ZN(new_n869));
  INV_X1    g683(.A(new_n690), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n497), .A3(new_n870), .A4(new_n865), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(KEYINPUT110), .A3(new_n659), .A4(new_n701), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n856), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n756), .A2(new_n766), .A3(new_n778), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n763), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n689), .A2(new_n691), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n713), .A2(new_n498), .A3(new_n754), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n676), .A2(new_n310), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n879), .A2(new_n881), .B1(new_n777), .B2(new_n775), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n882), .A3(KEYINPUT115), .A4(new_n766), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n794), .A2(new_n714), .A3(new_n598), .A4(new_n708), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n776), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n733), .B2(new_n729), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n716), .A2(new_n887), .A3(new_n747), .A4(new_n783), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT52), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n790), .A2(new_n781), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n715), .A2(new_n712), .B1(new_n890), .B2(new_n780), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n892), .A3(new_n747), .A4(new_n887), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n874), .A2(new_n884), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n868), .A2(new_n872), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n756), .A2(new_n766), .A3(new_n778), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n855), .A2(new_n897), .A3(new_n798), .A4(new_n880), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT111), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT111), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n876), .A2(new_n763), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n856), .A2(new_n873), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT112), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n889), .B2(new_n893), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n889), .A2(new_n893), .A3(new_n903), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n899), .B(new_n902), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n907));
  AOI211_X1 g721(.A(KEYINPUT54), .B(new_n895), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT114), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n899), .A2(new_n902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n905), .A2(new_n904), .ZN(new_n912));
  INV_X1    g726(.A(new_n907), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n899), .A2(new_n902), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n894), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n909), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n908), .B1(new_n918), .B2(KEYINPUT54), .ZN(new_n919));
  INV_X1    g733(.A(new_n817), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n792), .A2(new_n754), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n371), .A3(new_n782), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n371), .A3(new_n497), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n734), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n704), .A3(new_n745), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n817), .A2(new_n370), .A3(new_n773), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n682), .B1(KEYINPUT117), .B2(KEYINPUT50), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n754), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n720), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n922), .B(new_n925), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT51), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n846), .A2(KEYINPUT116), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n846), .A2(KEYINPUT116), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n599), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n832), .A2(new_n833), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT118), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n832), .A2(new_n940), .A3(new_n833), .A4(new_n937), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n926), .A2(new_n786), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n934), .A2(new_n943), .A3(KEYINPUT119), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT119), .B1(new_n934), .B2(new_n943), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n920), .A2(new_n371), .A3(new_n921), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT48), .ZN(new_n948));
  INV_X1    g762(.A(new_n597), .ZN(new_n949));
  OR4_X1    g763(.A1(KEYINPUT120), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n926), .A2(new_n780), .ZN(new_n951));
  INV_X1    g765(.A(G952), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n745), .A2(new_n704), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n952), .B(G953), .C1(new_n924), .C2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n947), .B2(new_n949), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n950), .A2(new_n951), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n938), .A2(new_n942), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n958), .A2(new_n932), .A3(new_n931), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(new_n933), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n919), .A2(new_n946), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(G952), .A2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n851), .B1(new_n961), .B2(new_n962), .ZN(G75));
  NAND2_X1  g777(.A1(new_n952), .A2(G953), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT121), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT56), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n905), .A2(new_n904), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n907), .B1(new_n916), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n895), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(G902), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n972), .B2(new_n306), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n253), .A2(new_n289), .A3(new_n290), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n288), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT55), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n973), .A2(new_n976), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n966), .B1(new_n977), .B2(new_n978), .ZN(G51));
  XNOR2_X1  g793(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n653), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT54), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n969), .B2(new_n970), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n908), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n752), .B2(new_n751), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n972), .A2(new_n804), .A3(new_n806), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n966), .B1(new_n985), .B2(new_n986), .ZN(G54));
  NAND2_X1  g801(.A1(KEYINPUT58), .A2(G475), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n972), .A2(new_n441), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n441), .B1(new_n972), .B2(new_n988), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n966), .B1(new_n989), .B2(new_n990), .ZN(G60));
  NAND2_X1  g805(.A1(G478), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT59), .Z(new_n993));
  NOR2_X1   g807(.A1(new_n672), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n908), .B2(new_n983), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT123), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT123), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n997), .B(new_n994), .C1(new_n908), .C2(new_n983), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n672), .B1(new_n919), .B2(new_n993), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n999), .A2(new_n965), .A3(new_n1000), .ZN(G63));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G217), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT124), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT60), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n971), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n696), .A2(new_n697), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT125), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n965), .B1(new_n1006), .B2(new_n495), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1002), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1006), .A2(new_n495), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1013), .A2(KEYINPUT61), .A3(new_n1009), .A4(new_n965), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(G66));
  OAI21_X1  g829(.A(G953), .B1(new_n285), .B2(new_n374), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n873), .A2(new_n901), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(G953), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n974), .B1(G898), .B2(new_n369), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G69));
  AOI21_X1  g834(.A(new_n369), .B1(G227), .B2(G900), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n558), .A2(new_n560), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT126), .Z(new_n1024));
  NAND2_X1  g838(.A1(new_n401), .A2(new_n402), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n706), .B2(new_n369), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n827), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n811), .A2(new_n597), .A3(new_n777), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n891), .A2(new_n747), .ZN(new_n1031));
  AND4_X1   g845(.A1(new_n798), .A2(new_n1030), .A3(new_n800), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n838), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1028), .B1(new_n1033), .B2(G953), .ZN(new_n1034));
  INV_X1    g848(.A(new_n865), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n658), .A2(new_n735), .ZN(new_n1036));
  NOR4_X1   g850(.A1(new_n949), .A2(new_n1035), .A3(new_n1036), .A4(new_n792), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1029), .A2(KEYINPUT127), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n738), .A2(new_n1031), .ZN(new_n1040));
  OR2_X1    g854(.A1(new_n1040), .A2(KEYINPUT62), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(KEYINPUT62), .ZN(new_n1042));
  AOI22_X1  g856(.A1(new_n836), .A2(new_n837), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT127), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1044), .B1(new_n827), .B2(new_n1037), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1039), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1046), .A2(new_n369), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1022), .B(new_n1034), .C1(new_n1047), .C2(new_n1026), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1026), .B1(new_n1046), .B2(new_n369), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1034), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1021), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1048), .A2(new_n1051), .ZN(G72));
  INV_X1    g866(.A(new_n726), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1039), .A2(new_n1043), .A3(new_n1017), .A4(new_n1045), .ZN(new_n1054));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  AOI21_X1  g870(.A(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n725), .A2(new_n503), .ZN(new_n1058));
  AND4_X1   g872(.A1(new_n1053), .A2(new_n918), .A3(new_n1058), .A4(new_n1056), .ZN(new_n1059));
  NAND4_X1  g873(.A1(new_n838), .A2(new_n1029), .A3(new_n1017), .A4(new_n1032), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1058), .B1(new_n1060), .B2(new_n1056), .ZN(new_n1061));
  NOR4_X1   g875(.A1(new_n1057), .A2(new_n1059), .A3(new_n966), .A4(new_n1061), .ZN(G57));
endmodule


