//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n448, new_n452,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g024(.A(G452), .Z(G391));
  AND2_X1   g025(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g028(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT2), .Z(new_n457));
  NAND4_X1  g032(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n470), .A2(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(new_n466), .B2(G136), .ZN(new_n477));
  INV_X1    g052(.A(new_n463), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n464), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n479), .A2(new_n480), .A3(G124), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n479), .B2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NOR2_X1   g059(.A1(new_n464), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n463), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n463), .A2(KEYINPUT71), .A3(new_n488), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n464), .A2(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n463), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n463), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n504), .B2(new_n505), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(G88), .B1(new_n508), .B2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(new_n503), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n509), .B1(new_n510), .B2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(G89), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(G51), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n522), .A2(new_n529), .ZN(G168));
  OAI211_X1 g105(.A(G52), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n516), .A2(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(G90), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G64), .B1(new_n515), .B2(new_n516), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n510), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  XNOR2_X1  g113(.A(KEYINPUT6), .B(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G43), .A3(G543), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  OAI21_X1  g117(.A(G56), .B1(new_n515), .B2(new_n516), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n510), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  INV_X1    g126(.A(new_n508), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n508), .A2(new_n555), .A3(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n532), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n511), .A2(new_n539), .A3(KEYINPUT73), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(G91), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT74), .B(G65), .Z(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(new_n517), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n557), .A2(new_n561), .A3(new_n565), .ZN(G299));
  OAI21_X1  g141(.A(KEYINPUT75), .B1(new_n534), .B2(new_n537), .ZN(new_n567));
  INV_X1    g142(.A(G64), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n502), .B2(new_n503), .ZN(new_n569));
  INV_X1    g144(.A(new_n536), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT72), .B(G90), .Z(new_n573));
  NAND3_X1  g148(.A1(new_n573), .A2(new_n511), .A3(new_n539), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n571), .A2(new_n572), .A3(new_n574), .A4(new_n531), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G301));
  INV_X1    g152(.A(G89), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n504), .B2(new_n505), .ZN(new_n579));
  INV_X1    g154(.A(new_n521), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n511), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(new_n528), .A3(new_n527), .ZN(G286));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  INV_X1    g158(.A(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n552), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n508), .A2(KEYINPUT76), .A3(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n559), .A2(G87), .A3(new_n560), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n559), .A2(G86), .A3(new_n560), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n517), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n508), .A2(G48), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n510), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n508), .A2(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n532), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(KEYINPUT77), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n506), .A2(G85), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n600), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n603), .B2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT78), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT80), .B(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n508), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n559), .A2(G92), .A3(new_n560), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT79), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n559), .A2(new_n617), .A3(G92), .A4(new_n560), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n615), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n609), .B1(G868), .B2(new_n622), .ZN(G284));
  OAI21_X1  g198(.A(new_n609), .B1(G868), .B2(new_n622), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n463), .A2(new_n468), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n479), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n466), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n464), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT81), .Z(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT83), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n665), .A3(new_n667), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n666), .A2(new_n667), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n665), .A2(new_n667), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n677), .A2(new_n669), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n672), .B(new_n675), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n686), .A2(new_n688), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n684), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n689), .A3(new_n684), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n690), .B1(new_n689), .B2(new_n684), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(G23), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n705), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n705), .A2(G6), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G305), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  AOI22_X1  g292(.A1(new_n711), .A2(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n714), .B(new_n718), .C1(new_n716), .C2(new_n717), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n721));
  MUX2_X1   g296(.A(G24), .B(G290), .S(G16), .Z(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT88), .Z(new_n723));
  INV_X1    g298(.A(G1986), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G25), .A2(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n479), .A2(G119), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n466), .A2(G131), .ZN(new_n728));
  OR2_X1    g303(.A1(G95), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT87), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n723), .B2(new_n724), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n720), .A2(new_n721), .A3(new_n725), .A4(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT36), .Z(new_n739));
  NAND2_X1  g314(.A1(G115), .A2(G2104), .ZN(new_n740));
  INV_X1    g315(.A(G127), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n478), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G2105), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G139), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n465), .ZN(new_n748));
  OAI21_X1  g323(.A(G29), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G33), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(new_n444), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT93), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT26), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n479), .B2(G129), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n466), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G32), .B(new_n760), .S(G29), .Z(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT95), .Z(new_n762));
  AOI21_X1  g337(.A(new_n754), .B1(new_n755), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n705), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n626), .B2(new_n705), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT101), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G1956), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n763), .B(new_n769), .C1(new_n755), .C2(new_n762), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G35), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G162), .B2(G29), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2090), .ZN(new_n775));
  AND2_X1   g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NOR2_X1   g351(.A1(KEYINPUT24), .A2(G34), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n750), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT94), .Z(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n472), .B2(new_n750), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n752), .A2(new_n444), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  NOR2_X1   g359(.A1(G171), .A2(new_n705), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G5), .B2(new_n705), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n750), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n750), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n789), .A2(G2078), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(G2078), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT96), .B1(new_n644), .B2(new_n750), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT97), .B(G28), .Z(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(new_n750), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n792), .B(new_n793), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n644), .A2(KEYINPUT96), .A3(new_n750), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n790), .A2(new_n791), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n786), .A2(new_n784), .B1(new_n780), .B2(new_n781), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n705), .A2(G21), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G168), .B2(new_n705), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1966), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n775), .A2(new_n787), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n770), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G4), .A2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT89), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n621), .B2(new_n705), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT90), .B(G1348), .Z(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n705), .A2(G19), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n546), .B2(new_n705), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1341), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n750), .A2(G26), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT91), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT28), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n479), .A2(G128), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n466), .A2(G140), .ZN(new_n821));
  OR2_X1    g396(.A1(G104), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(new_n750), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2067), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n812), .A2(new_n813), .A3(new_n816), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  OR3_X1    g405(.A1(new_n774), .A2(new_n830), .A3(G2090), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n768), .A2(G1956), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n830), .B1(new_n774), .B2(G2090), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n807), .A2(new_n829), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n770), .A2(new_n834), .A3(new_n806), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n840), .A2(KEYINPUT102), .A3(new_n829), .A4(new_n836), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n739), .B1(new_n839), .B2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n739), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n508), .A2(G55), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n511), .A2(new_n539), .A3(G93), .ZN(new_n848));
  OAI21_X1  g423(.A(G67), .B1(new_n515), .B2(new_n516), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n510), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n847), .B(new_n848), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n854), .A2(KEYINPUT103), .A3(new_n510), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n846), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT103), .B1(new_n854), .B2(new_n510), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n847), .A2(new_n848), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n852), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT105), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n622), .A2(G559), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT106), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  INV_X1    g441(.A(new_n546), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n856), .A2(new_n867), .A3(new_n860), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n546), .B1(new_n853), .B2(new_n855), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(KEYINPUT104), .A3(new_n546), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n865), .B(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n869), .A2(new_n870), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT104), .B1(new_n872), .B2(new_n546), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n868), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n875), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G860), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n875), .B2(new_n881), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n863), .B1(new_n885), .B2(new_n886), .ZN(G145));
  NOR2_X1   g462(.A1(new_n743), .A2(new_n748), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n760), .Z(new_n889));
  AOI22_X1  g464(.A1(G130), .A2(new_n479), .B1(new_n466), .B2(G142), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n464), .A2(G118), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n467), .B1(new_n891), .B2(KEYINPUT108), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT108), .B1(G106), .B2(G2105), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(new_n636), .Z(new_n897));
  XOR2_X1   g472(.A(new_n889), .B(new_n897), .Z(new_n898));
  INV_X1    g473(.A(new_n492), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT71), .B1(new_n463), .B2(new_n488), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n899), .A2(new_n900), .B1(new_n485), .B2(new_n486), .ZN(new_n901));
  INV_X1    g476(.A(new_n498), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n497), .B1(new_n463), .B2(new_n494), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT107), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n496), .A2(new_n905), .A3(new_n498), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n825), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n731), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n889), .B(new_n897), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n644), .B(new_n472), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(G162), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n916), .A3(new_n913), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n918), .A2(new_n923), .A3(new_n919), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n512), .A2(new_n510), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n508), .A2(G50), .ZN(new_n929));
  INV_X1    g504(.A(G88), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(new_n532), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n509), .B(KEYINPUT110), .C1(new_n510), .C2(new_n512), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n710), .ZN(new_n935));
  NAND3_X1  g510(.A1(G288), .A2(new_n932), .A3(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G305), .ZN(new_n938));
  NAND2_X1  g513(.A1(G290), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(G305), .B(new_n599), .C1(new_n603), .C2(new_n606), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n935), .A2(new_n939), .A3(new_n940), .A4(new_n936), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT42), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n631), .B(new_n880), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n615), .A2(new_n618), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT10), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n626), .B1(new_n951), .B2(new_n613), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n626), .B(new_n613), .C1(new_n619), .C2(new_n620), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n947), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n952), .B2(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n621), .A2(G299), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(KEYINPUT41), .A3(new_n953), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n947), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n946), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n946), .B1(new_n957), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G868), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n861), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(G295));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n966), .A2(new_n970), .A3(new_n968), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n966), .B2(new_n968), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(G331));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n974));
  NOR2_X1   g549(.A1(KEYINPUT43), .A2(G37), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n567), .A2(new_n575), .A3(G168), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(G171), .B2(G286), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n567), .A2(new_n575), .A3(new_n977), .A4(G168), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n880), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n567), .A2(G168), .A3(new_n575), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n571), .A2(new_n531), .A3(new_n574), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT112), .B1(new_n984), .B2(G168), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n980), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n874), .A2(new_n986), .A3(new_n868), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n959), .A2(new_n961), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n982), .A2(new_n960), .A3(new_n987), .A4(new_n953), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n944), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n975), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n959), .A2(new_n988), .A3(new_n961), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n944), .B1(new_n993), .B2(new_n990), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n974), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n919), .B1(new_n989), .B2(new_n991), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT43), .B1(new_n996), .B2(new_n994), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n990), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n942), .A2(new_n943), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n975), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n874), .A2(new_n986), .A3(new_n868), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n986), .B1(new_n868), .B2(new_n874), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n999), .B1(new_n1004), .B2(new_n955), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n1005), .B2(new_n993), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1006), .A3(KEYINPUT113), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n995), .A2(new_n997), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT114), .B1(new_n996), .B2(new_n994), .ZN(new_n1011));
  AOI21_X1  g586(.A(G37), .B1(new_n1005), .B2(new_n993), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1000), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(KEYINPUT43), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1009), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1010), .A2(new_n1017), .A3(KEYINPUT115), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(G397));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n907), .B2(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n469), .A2(new_n471), .A3(G40), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n731), .B(new_n734), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1027), .A2(KEYINPUT116), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(KEYINPUT116), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n824), .A2(G2067), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n824), .A2(G2067), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1996), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n760), .B(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(G290), .B(G1986), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1026), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n904), .A2(new_n906), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n493), .ZN(new_n1041));
  INV_X1    g616(.A(G1384), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1025), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1023), .A2(G1384), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(G164), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1039), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT121), .B(new_n1039), .C1(new_n1043), .C2(new_n1047), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n907), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1384), .B1(new_n493), .B2(new_n499), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1044), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n781), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1051), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT118), .B(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G168), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1038), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1038), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1060), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1058), .A2(new_n1067), .A3(new_n1061), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1063), .A2(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  OAI221_X1 g648(.A(new_n1073), .B1(new_n1069), .B2(new_n1070), .C1(new_n1063), .C2(new_n1066), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G303), .A2(G8), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT55), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1971), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1044), .B1(new_n907), .B2(new_n1046), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1053), .A2(KEYINPUT45), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT117), .B(new_n1078), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n500), .A2(new_n1042), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1025), .B1(new_n1082), .B2(KEYINPUT50), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1084), .B2(KEYINPUT50), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1081), .B1(new_n1085), .B2(G2090), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1025), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1023), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1971), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(KEYINPUT117), .ZN(new_n1090));
  OAI211_X1 g665(.A(G8), .B(new_n1077), .C1(new_n1086), .C2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1054), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1044), .B1(new_n1082), .B2(KEYINPUT50), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(G2090), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1065), .B1(new_n1094), .B2(new_n1089), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1076), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1044), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n710), .A2(G1976), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1065), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT52), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(KEYINPUT119), .A3(KEYINPUT52), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n710), .B2(G1976), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1981), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n591), .A2(new_n1108), .A3(new_n595), .A4(new_n596), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT120), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n506), .A2(G86), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n595), .A2(new_n596), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G1981), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT49), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1097), .A2(new_n1065), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1110), .A2(KEYINPUT49), .A3(new_n1113), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1107), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1091), .A2(new_n1096), .A3(new_n1104), .A4(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1087), .A2(new_n445), .A3(new_n1088), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n784), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1025), .B1(new_n500), .B2(new_n1045), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1024), .A2(KEYINPUT53), .A3(new_n1124), .A4(new_n445), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n576), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1119), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1072), .A2(new_n1074), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT54), .B1(new_n1126), .B2(new_n576), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n784), .A2(new_n1085), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1087), .A2(new_n1024), .A3(KEYINPUT53), .A4(new_n445), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n984), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1122), .A2(new_n1123), .A3(G301), .A4(new_n1132), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT54), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1134), .A2(new_n1119), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1956), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1087), .A2(new_n1088), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(G299), .B(KEYINPUT57), .Z(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1056), .A2(G1348), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1097), .A2(G2067), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1148), .B2(new_n621), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1139), .A2(new_n1143), .A3(new_n1141), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1153));
  OAI221_X1 g728(.A(KEYINPUT60), .B1(G2067), .B2(new_n1097), .C1(new_n1056), .C2(G1348), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n622), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1150), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1143), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1145), .A2(new_n1150), .A3(KEYINPUT61), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1087), .A2(new_n1033), .A3(new_n1088), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1097), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT58), .B(G1341), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n546), .ZN(new_n1166));
  NAND2_X1  g741(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1165), .A2(KEYINPUT123), .A3(KEYINPUT59), .A4(new_n546), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1168), .B(new_n1169), .C1(new_n622), .C2(new_n1154), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1151), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1137), .A2(new_n1171), .A3(new_n1071), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1118), .A2(new_n1104), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1110), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1175));
  NOR2_X1   g750(.A1(G288), .A2(G1976), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1173), .A2(new_n1091), .B1(new_n1177), .B2(new_n1115), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1058), .A2(G168), .A3(new_n1065), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1119), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1118), .A2(new_n1104), .A3(KEYINPUT63), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1180), .ZN(new_n1183));
  OAI21_X1  g758(.A(G8), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(KEYINPUT122), .A3(new_n1076), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1076), .A2(KEYINPUT122), .ZN(new_n1186));
  OAI211_X1 g761(.A(G8), .B(new_n1186), .C1(new_n1086), .C2(new_n1090), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1178), .B1(new_n1181), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1172), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1037), .B1(new_n1129), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n732), .A2(new_n734), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1030), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1026), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1026), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1196), .A2(G1986), .A3(G290), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT126), .Z(new_n1198));
  INV_X1    g773(.A(KEYINPUT48), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1035), .A2(new_n1026), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1195), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT46), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(new_n1196), .B2(G1996), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1032), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1026), .B1(new_n1206), .B2(new_n760), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1026), .A2(KEYINPUT46), .A3(new_n1033), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT47), .Z(new_n1210));
  AND2_X1   g785(.A1(new_n1210), .A2(KEYINPUT125), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1210), .A2(KEYINPUT125), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1203), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1191), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g789(.A(G319), .B1(new_n662), .B2(new_n663), .ZN(new_n1216));
  OR3_X1    g790(.A1(G227), .A2(KEYINPUT127), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g791(.A(KEYINPUT127), .B1(G227), .B2(new_n1216), .ZN(new_n1218));
  AND3_X1   g792(.A1(new_n1217), .A2(new_n703), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n1219), .A2(new_n925), .A3(new_n1008), .ZN(G225));
  INV_X1    g794(.A(G225), .ZN(G308));
endmodule


