//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G1gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n208), .B(KEYINPUT91), .C1(new_n209), .C2(G1gat), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n213), .A2(KEYINPUT92), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G15gat), .B(G22gat), .Z(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n219), .B(new_n210), .C1(new_n212), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G8gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT89), .B1(new_n224), .B2(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT15), .ZN(new_n228));
  INV_X1    g027(.A(G43gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G50gat), .ZN(new_n230));
  INV_X1    g029(.A(G50gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G43gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n227), .B(new_n228), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT88), .B(G29gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G36gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT14), .ZN(new_n238));
  INV_X1    g037(.A(G29gat), .ZN(new_n239));
  INV_X1    g038(.A(G36gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT90), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n237), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(G29gat), .A2(G36gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT90), .B1(new_n244), .B2(new_n238), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n236), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n225), .B1(new_n234), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n225), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n241), .A2(KEYINPUT87), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n237), .B1(new_n241), .B2(KEYINPUT87), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n248), .B(new_n236), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n247), .A2(KEYINPUT17), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT17), .B1(new_n247), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n223), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G229gat), .A2(G233gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n251), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n216), .A2(new_n222), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n207), .B1(new_n263), .B2(KEYINPUT95), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n223), .A2(new_n256), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT94), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n255), .B(KEYINPUT13), .Z(new_n268));
  NAND3_X1  g067(.A1(new_n223), .A2(KEYINPUT94), .A3(new_n256), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n254), .A2(KEYINPUT18), .A3(new_n255), .A4(new_n259), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n264), .A2(new_n272), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT96), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n263), .A2(KEYINPUT95), .ZN(new_n277));
  INV_X1    g076(.A(new_n207), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n263), .A2(new_n270), .A3(new_n271), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n272), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT96), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  INV_X1    g085(.A(G113gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n288));
  INV_X1    g087(.A(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT66), .B1(new_n287), .B2(G120gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n285), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G127gat), .B(G134gat), .Z(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(KEYINPUT1), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G141gat), .ZN(new_n306));
  INV_X1    g105(.A(G141gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n303), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n304), .B1(new_n303), .B2(new_n309), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT72), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(G155gat), .B2(G162gat), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n307), .A2(G148gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n305), .A2(G141gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n298), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n319), .A3(new_n302), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n297), .A2(new_n312), .A3(KEYINPUT4), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  AND2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n298), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G141gat), .B(G148gat), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT73), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n303), .A2(new_n304), .A3(new_n309), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n320), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n293), .A2(new_n296), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n322), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(new_n312), .B2(new_n320), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n320), .A2(new_n327), .A3(new_n332), .A4(new_n328), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n330), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n321), .B(new_n331), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT75), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n321), .A2(new_n331), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(new_n330), .A3(new_n334), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n339), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n297), .A2(new_n312), .A3(new_n320), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n330), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n351), .A3(new_n330), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n338), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n322), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n353), .B(KEYINPUT5), .C1(new_n336), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT81), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n355), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n355), .A3(new_n361), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(KEYINPUT22), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G211gat), .B(G218gat), .Z(new_n375));
  OR2_X1    g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n375), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G190gat), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT28), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT27), .B(G183gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT28), .A3(new_n381), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390));
  INV_X1    g189(.A(G169gat), .ZN(new_n391));
  INV_X1    g190(.A(G176gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399));
  AND2_X1   g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(KEYINPUT24), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT24), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT25), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT23), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n405), .A2(G169gat), .A3(G176gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n392), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n394), .A2(KEYINPUT23), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n389), .A2(new_n398), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n397), .A2(KEYINPUT64), .A3(new_n402), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT64), .ZN(new_n412));
  OAI211_X1 g211(.A(G183gat), .B(G190gat), .C1(new_n412), .C2(KEYINPUT24), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n411), .B(new_n413), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n409), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT25), .ZN(new_n419));
  AOI211_X1 g218(.A(KEYINPUT29), .B(new_n380), .C1(new_n410), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n410), .A2(new_n380), .A3(new_n419), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n378), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT71), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n378), .B(KEYINPUT70), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n389), .A2(new_n398), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n409), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n379), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n430), .A3(new_n421), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT71), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n378), .ZN(new_n434));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435));
  INV_X1    g234(.A(G64gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n437), .B(G92gat), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n424), .A2(new_n431), .A3(new_n434), .A4(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n433), .B1(new_n432), .B2(new_n378), .ZN(new_n442));
  INV_X1    g241(.A(new_n378), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT71), .B(new_n443), .C1(new_n430), .C2(new_n421), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT70), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n378), .B(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n432), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT37), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n439), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n432), .A2(new_n443), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n425), .B2(new_n432), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT38), .B1(new_n452), .B2(KEYINPUT37), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n441), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n356), .A2(new_n362), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n369), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n450), .B1(new_n449), .B2(new_n448), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT38), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n369), .A2(new_n454), .A3(KEYINPUT82), .A4(new_n457), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n334), .A2(new_n429), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n333), .B1(new_n425), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G228gat), .ZN(new_n467));
  INV_X1    g266(.A(G233gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n376), .B2(new_n377), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n329), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n471), .A2(KEYINPUT77), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n332), .B1(new_n471), .B2(KEYINPUT77), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n329), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n443), .A2(new_n465), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(G22gat), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n477), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n470), .ZN(new_n481));
  INV_X1    g280(.A(G22gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n480), .A2(new_n470), .B1(new_n466), .B2(new_n472), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT78), .B1(new_n486), .B2(new_n482), .ZN(new_n487));
  XNOR2_X1  g286(.A(G78gat), .B(G106gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT31), .B(G50gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n485), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n479), .A2(new_n484), .A3(KEYINPUT78), .A4(new_n490), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n424), .A2(new_n431), .A3(new_n434), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n438), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT30), .A3(new_n440), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n448), .A2(new_n498), .A3(new_n439), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n497), .A2(KEYINPUT79), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT79), .B1(new_n497), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n336), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT80), .B1(new_n503), .B2(new_n337), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n336), .A2(new_n505), .A3(new_n338), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n362), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n350), .A2(new_n352), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n510), .B2(new_n337), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n504), .A2(new_n511), .A3(new_n506), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT40), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n515), .A3(new_n512), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n361), .B1(new_n356), .B2(KEYINPUT81), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n514), .A2(new_n516), .B1(new_n364), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n494), .B1(new_n502), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n464), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT76), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n366), .A2(new_n367), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n456), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n368), .A2(KEYINPUT76), .A3(new_n455), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n457), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n497), .A2(new_n499), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n494), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n428), .B2(new_n330), .ZN(new_n531));
  NAND2_X1  g330(.A1(G227gat), .A2(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n428), .A2(new_n330), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n410), .A2(KEYINPUT67), .A3(new_n297), .A4(new_n419), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT34), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT32), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(new_n532), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT33), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G43gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G71gat), .B(G99gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n536), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(new_n539), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT32), .ZN(new_n551));
  INV_X1    g350(.A(new_n541), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n544), .ZN(new_n553));
  INV_X1    g352(.A(new_n536), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT69), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n549), .A2(new_n555), .A3(KEYINPUT68), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n536), .C1(new_n547), .C2(new_n548), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n557), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n464), .A2(new_n519), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n521), .A2(new_n529), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n565), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n492), .A2(new_n493), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n526), .A3(new_n527), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT85), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n369), .A2(new_n457), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n494), .A2(new_n556), .ZN(new_n580));
  INV_X1    g379(.A(new_n502), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n582));
  AND4_X1   g381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n284), .B1(new_n570), .B2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G71gat), .B(G78gat), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n436), .A2(G57gat), .ZN(new_n589));
  INV_X1    g388(.A(G57gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G64gat), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT97), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT97), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n588), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n591), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n597), .A2(new_n588), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n223), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT100), .ZN(new_n604));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT99), .B(KEYINPUT21), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n604), .B(new_n605), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n611), .A2(new_n614), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT101), .Z(new_n624));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n381), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n372), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n624), .A2(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n256), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n247), .A2(KEYINPUT17), .A3(new_n251), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G85gat), .ZN(new_n638));
  AND2_X1   g437(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G99gat), .ZN(new_n642));
  INV_X1    g441(.A(G106gat), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT8), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G99gat), .B(G106gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n637), .A2(new_n641), .A3(new_n646), .A4(new_n644), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n630), .B1(new_n634), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n257), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n651), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n629), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n628), .B(G218gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n656), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n650), .B1(new_n598), .B2(new_n600), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n599), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n595), .A2(KEYINPUT98), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n595), .A2(KEYINPUT98), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT97), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n587), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n597), .A2(new_n588), .A3(new_n599), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n649), .A4(new_n648), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n664), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n654), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n673), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(G230gat), .A3(G233gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT104), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n289), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n679), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n678), .B(KEYINPUT105), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n677), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n685), .B1(new_n689), .B2(new_n681), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n622), .A2(new_n663), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT106), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n622), .A2(new_n695), .A3(new_n663), .A4(new_n692), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT107), .B1(new_n586), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n586), .A2(KEYINPUT107), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n526), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g503(.A1(new_n209), .A2(new_n214), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n701), .A2(new_n502), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n209), .A2(new_n214), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n701), .ZN(new_n710));
  OAI21_X1  g509(.A(G8gat), .B1(new_n710), .B2(new_n581), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(G1325gat));
  INV_X1    g512(.A(new_n556), .ZN(new_n714));
  AOI21_X1  g513(.A(G15gat), .B1(new_n701), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n710), .A2(new_n567), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n494), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  INV_X1    g520(.A(new_n663), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n464), .A2(new_n519), .A3(new_n568), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n568), .B1(new_n464), .B2(new_n519), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n529), .B1(new_n562), .B2(new_n566), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n721), .B(new_n722), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n570), .A2(new_n585), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n731), .A2(new_n721), .A3(KEYINPUT44), .A4(new_n722), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n281), .A2(new_n282), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n622), .A2(new_n691), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n235), .B1(new_n735), .B2(new_n526), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n722), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n526), .A2(new_n235), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n586), .A2(new_n739), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1328gat));
  AND3_X1   g545(.A1(new_n586), .A2(new_n739), .A3(new_n740), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n240), .A3(new_n502), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT46), .Z(new_n749));
  OAI21_X1  g548(.A(G36gat), .B1(new_n735), .B2(new_n581), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1329gat));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  OAI21_X1  g551(.A(G43gat), .B1(new_n735), .B2(new_n567), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n747), .A2(new_n229), .A3(new_n714), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1330gat));
  AOI21_X1  g556(.A(G50gat), .B1(new_n747), .B2(new_n494), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n735), .A2(new_n231), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n494), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1331gat));
  INV_X1    g561(.A(new_n733), .ZN(new_n763));
  INV_X1    g562(.A(new_n622), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n722), .A3(new_n692), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n731), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n526), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n590), .ZN(G1332gat));
  AOI21_X1  g567(.A(new_n581), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT112), .Z(new_n770));
  NOR2_X1   g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT113), .Z(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1333gat));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  INV_X1    g574(.A(G71gat), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n766), .A2(new_n776), .A3(new_n567), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n766), .B2(new_n556), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n775), .A3(new_n778), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n780), .A2(KEYINPUT50), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT50), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n766), .A2(new_n572), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(G78gat), .Z(G1335gat));
  AND2_X1   g585(.A1(new_n730), .A2(new_n732), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n622), .A2(new_n733), .A3(new_n692), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(new_n638), .A3(new_n526), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n622), .A2(new_n733), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n722), .B(new_n791), .C1(new_n726), .C2(new_n727), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n722), .A4(new_n791), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n692), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n702), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n790), .A2(new_n797), .ZN(G1336gat));
  NOR2_X1   g597(.A1(new_n581), .A2(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n730), .A2(new_n732), .A3(new_n502), .A4(new_n788), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n639), .A2(new_n640), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n799), .A2(new_n691), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n794), .B2(new_n795), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT115), .B1(new_n792), .B2(new_n793), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n803), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n806), .B1(new_n813), .B2(KEYINPUT52), .ZN(new_n814));
  AOI211_X1 g613(.A(KEYINPUT116), .B(new_n804), .C1(new_n812), .C2(new_n803), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n805), .B1(new_n814), .B2(new_n815), .ZN(G1337gat));
  OAI21_X1  g615(.A(G99gat), .B1(new_n789), .B2(new_n567), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n796), .A2(new_n642), .A3(new_n714), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1338gat));
  NAND3_X1  g618(.A1(new_n787), .A2(new_n494), .A3(new_n788), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n796), .A2(new_n643), .A3(new_n494), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n810), .A2(new_n811), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n572), .A2(G106gat), .A3(new_n692), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n825), .A2(new_n826), .B1(new_n820), .B2(G106gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n822), .ZN(G1339gat));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n677), .A2(new_n831), .A3(new_n688), .ZN(new_n832));
  INV_X1    g631(.A(new_n685), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n830), .A3(new_n833), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n679), .B(KEYINPUT54), .C1(new_n677), .C2(new_n688), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n832), .A2(new_n830), .A3(new_n833), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT55), .B(new_n838), .C1(new_n841), .C2(new_n834), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(KEYINPUT118), .A3(new_n686), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT118), .B1(new_n842), .B2(new_n686), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n840), .B(new_n733), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n280), .A2(new_n207), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n255), .B1(new_n254), .B2(new_n259), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n206), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n846), .A2(new_n691), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n722), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n839), .A2(new_n663), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n846), .A2(new_n849), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n853), .B(new_n854), .C1(new_n844), .C2(new_n843), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n829), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n686), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n842), .A2(KEYINPUT118), .A3(new_n686), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n839), .B1(new_n281), .B2(new_n282), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n850), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT119), .B(new_n855), .C1(new_n864), .C2(new_n722), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n764), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n622), .A2(new_n763), .A3(new_n663), .A4(new_n692), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n580), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n502), .A2(new_n526), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n284), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n868), .A2(new_n572), .A3(new_n571), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n870), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n287), .A3(new_n733), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n877), .ZN(G1340gat));
  OAI21_X1  g677(.A(G120gat), .B1(new_n872), .B2(new_n692), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n289), .A3(new_n691), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n871), .A2(G127gat), .A3(new_n622), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT120), .Z(new_n883));
  AOI21_X1  g682(.A(G127gat), .B1(new_n876), .B2(new_n622), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(G1342gat));
  INV_X1    g684(.A(G134gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n502), .A2(new_n663), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT121), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n874), .A2(new_n886), .A3(new_n702), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT56), .Z(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n872), .B2(new_n663), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1343gat));
  AOI211_X1 g691(.A(KEYINPUT57), .B(new_n572), .C1(new_n866), .C2(new_n867), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n567), .A2(new_n870), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n858), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n840), .B(new_n896), .C1(new_n276), .C2(new_n283), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n722), .B1(new_n897), .B2(new_n851), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n764), .B1(new_n898), .B2(new_n856), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n572), .B1(new_n899), .B2(new_n867), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n895), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n893), .A2(new_n902), .A3(KEYINPUT122), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n275), .B1(new_n273), .B2(new_n274), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n281), .A2(KEYINPUT96), .A3(new_n282), .ZN(new_n906));
  AOI211_X1 g705(.A(new_n839), .B(new_n858), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n663), .B1(new_n907), .B2(new_n850), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n622), .B1(new_n908), .B2(new_n855), .ZN(new_n909));
  INV_X1    g708(.A(new_n867), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n494), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n894), .B1(new_n911), .B2(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n868), .A2(new_n901), .A3(new_n494), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n733), .B1(new_n903), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(KEYINPUT123), .A3(G141gat), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT122), .B1(new_n893), .B2(new_n902), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n904), .A3(new_n913), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n763), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(new_n307), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n868), .A2(new_n494), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n894), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n284), .A2(G141gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n916), .A2(new_n921), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT58), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n913), .ZN(new_n930));
  OAI21_X1  g729(.A(G141gat), .B1(new_n930), .B2(new_n284), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(new_n925), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n929), .A2(new_n935), .ZN(G1344gat));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n937));
  AOI211_X1 g736(.A(new_n937), .B(G148gat), .C1(new_n923), .C2(new_n691), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n903), .A2(new_n914), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n937), .B1(new_n939), .B2(new_n692), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n694), .A2(new_n284), .A3(new_n696), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT57), .B1(new_n941), .B2(new_n899), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n922), .A2(KEYINPUT57), .B1(new_n942), .B2(new_n494), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n691), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n895), .A2(KEYINPUT59), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n938), .B1(new_n946), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g746(.A(G155gat), .B1(new_n923), .B2(new_n622), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n939), .A2(new_n764), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g749(.A(G162gat), .B1(new_n939), .B2(new_n663), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n888), .A2(new_n300), .A3(new_n702), .A4(new_n567), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n922), .B2(new_n952), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n581), .A2(new_n702), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n869), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G169gat), .B1(new_n956), .B2(new_n284), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n874), .A2(new_n954), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n391), .A3(new_n733), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1348gat));
  AOI21_X1  g759(.A(G176gat), .B1(new_n958), .B2(new_n691), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n956), .A2(new_n692), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(G176gat), .ZN(G1349gat));
  NAND2_X1  g762(.A1(new_n955), .A2(new_n622), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n622), .A2(new_n387), .ZN(new_n965));
  AOI22_X1  g764(.A1(new_n964), .A2(G183gat), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n381), .B1(new_n955), .B2(new_n722), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(KEYINPUT126), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(KEYINPUT126), .B2(new_n969), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n958), .A2(new_n381), .A3(new_n722), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n969), .A2(KEYINPUT126), .A3(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n941), .A2(new_n899), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n901), .A3(new_n494), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n567), .A2(new_n954), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n572), .B1(new_n866), .B2(new_n867), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n976), .B(new_n978), .C1(new_n979), .C2(new_n901), .ZN(new_n980));
  OAI21_X1  g779(.A(G197gat), .B1(new_n980), .B2(new_n284), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n922), .A2(new_n977), .ZN(new_n982));
  INV_X1    g781(.A(G197gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n983), .A3(new_n733), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n981), .A2(new_n984), .ZN(G1352gat));
  NOR4_X1   g784(.A1(new_n922), .A2(G204gat), .A3(new_n692), .A4(new_n977), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  OAI21_X1  g786(.A(G204gat), .B1(new_n944), .B2(new_n977), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1353gat));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(new_n980), .B2(new_n764), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n943), .A2(KEYINPUT127), .A3(new_n622), .A4(new_n978), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n991), .A2(G211gat), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n982), .A2(new_n371), .A3(new_n622), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n980), .B2(new_n663), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n372), .A3(new_n722), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1355gat));
endmodule


