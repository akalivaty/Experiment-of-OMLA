//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n212), .B(KEYINPUT25), .C1(G169gat), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G183gat), .B(G190gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(new_n219), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n224), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT65), .B(G169gat), .Z(new_n227));
  AND2_X1   g026(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .A4(new_n212), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n234), .A2(KEYINPUT26), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(KEYINPUT26), .ZN(new_n236));
  AOI211_X1 g035(.A(new_n218), .B(new_n235), .C1(new_n210), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n217), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(KEYINPUT66), .A2(KEYINPUT27), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT66), .A2(KEYINPUT27), .ZN(new_n245));
  OAI21_X1  g044(.A(G183gat), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n246), .B2(KEYINPUT67), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(G183gat), .C1(new_n244), .C2(new_n245), .ZN(new_n249));
  AOI221_X4 g048(.A(KEYINPUT68), .B1(KEYINPUT28), .B2(new_n241), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g051(.A(new_n243), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(KEYINPUT28), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n237), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n233), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT69), .B(new_n237), .C1(new_n250), .C2(new_n256), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n232), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n209), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n260), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT76), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT76), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(new_n260), .C1(new_n265), .C2(KEYINPUT29), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n260), .B1(new_n233), .B2(new_n257), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n268), .B1(new_n275), .B2(new_n209), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n209), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n273), .B1(new_n269), .B2(KEYINPUT76), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT77), .B1(new_n285), .B2(new_n268), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n278), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G85gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G141gat), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G148gat), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT79), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G155gat), .B(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT2), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n296), .B2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G120gat), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT1), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(G127gat), .A2(G134gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G127gat), .A2(G134gat), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT70), .B1(new_n309), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n310), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n308), .C1(new_n311), .C2(new_n312), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n303), .A2(new_n314), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n316), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n323), .A2(KEYINPUT82), .A3(new_n303), .A4(new_n314), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n325));
  INV_X1    g124(.A(new_n303), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n301), .B2(new_n302), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n296), .A2(new_n300), .ZN(new_n335));
  INV_X1    g134(.A(new_n297), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n317), .B1(new_n344), .B2(new_n308), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n334), .B(new_n340), .C1(new_n322), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT81), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n325), .A2(new_n348), .A3(new_n340), .A4(new_n334), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n321), .A2(new_n324), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n319), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n350), .A2(new_n352), .A3(new_n329), .A4(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n328), .A2(KEYINPUT83), .A3(new_n330), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n333), .A2(KEYINPUT5), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n321), .A2(new_n324), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT4), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  AOI211_X1 g162(.A(KEYINPUT5), .B(new_n330), .C1(new_n347), .C2(new_n349), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n351), .B1(new_n321), .B2(new_n324), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT84), .B1(new_n365), .B2(new_n361), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n291), .B1(new_n357), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n357), .A2(new_n367), .A3(new_n291), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n373), .A3(KEYINPUT6), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n368), .B2(KEYINPUT6), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n285), .A2(new_n268), .A3(new_n282), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT30), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n287), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n276), .B2(new_n281), .ZN(new_n382));
  NOR4_X1   g181(.A1(new_n285), .A2(KEYINPUT78), .A3(new_n268), .A4(new_n282), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT30), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n202), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n276), .A2(new_n281), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n378), .A2(new_n381), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n367), .ZN(new_n391));
  INV_X1    g190(.A(new_n291), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(KEYINPUT6), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT85), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n374), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n372), .B1(new_n378), .B2(KEYINPUT30), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n390), .A2(new_n396), .A3(KEYINPUT86), .A4(new_n287), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n340), .A2(new_n259), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n209), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n209), .A2(KEYINPUT29), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(new_n303), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(G228gat), .A3(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n339), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n326), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n406), .C1(KEYINPUT88), .C2(new_n399), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n399), .A2(KEYINPUT88), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  INV_X1    g211(.A(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G22gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n411), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n263), .A2(new_n264), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n233), .ZN(new_n418));
  INV_X1    g217(.A(new_n325), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G227gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n265), .A2(new_n325), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT32), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G15gat), .B(G43gat), .Z(new_n429));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n425), .B(KEYINPUT32), .C1(new_n427), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT74), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n424), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT72), .ZN(new_n440));
  INV_X1    g239(.A(new_n423), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n442), .A3(new_n424), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n423), .A2(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT73), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n439), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n444), .A2(KEYINPUT34), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n436), .A2(new_n438), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(KEYINPUT34), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n454), .A2(new_n437), .A3(new_n432), .A4(new_n434), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n416), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n385), .A2(new_n397), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n287), .A2(new_n379), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n384), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT35), .B1(new_n395), .B2(new_n372), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n460), .A2(new_n456), .A3(KEYINPUT90), .A4(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n458), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n385), .A2(new_n397), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n416), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n455), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n451), .A2(new_n455), .A3(new_n471), .A4(KEYINPUT36), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT37), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n281), .B1(new_n276), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n275), .A2(new_n283), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n261), .A2(new_n267), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n481), .B(KEYINPUT37), .C1(new_n283), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n278), .A2(KEYINPUT37), .A3(new_n286), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n485), .A2(new_n479), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n477), .B(new_n484), .C1(new_n486), .C2(new_n480), .ZN(new_n487));
  INV_X1    g286(.A(new_n416), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n363), .A2(new_n366), .A3(new_n350), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n330), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(KEYINPUT39), .C1(new_n330), .C2(new_n328), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT39), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n492), .A3(new_n330), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n493), .A2(new_n494), .A3(new_n291), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n493), .B2(new_n291), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT40), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n368), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n499), .B(new_n500), .C1(new_n384), .C2(new_n459), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n487), .A2(new_n488), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n469), .A2(new_n476), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n466), .A2(new_n467), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n467), .B1(new_n466), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  NOR2_X1   g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT14), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n510), .A2(KEYINPUT92), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n510), .B2(KEYINPUT92), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(KEYINPUT15), .B2(new_n507), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n510), .B(KEYINPUT93), .Z(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(G1gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(KEYINPUT16), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526));
  AOI211_X1 g325(.A(G8gat), .B(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(G8gat), .B1(new_n525), .B2(new_n522), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n527), .A2(new_n528), .B1(KEYINPUT94), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(KEYINPUT94), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n531), .B2(new_n518), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n531), .B(new_n518), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n534), .B(KEYINPUT13), .Z(new_n538));
  AOI22_X1  g337(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n534), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G197gat), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT11), .B(G169gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT12), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n539), .A2(new_n548), .A3(new_n540), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT96), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(KEYINPUT96), .A3(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n506), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G71gat), .B(G78gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT97), .Z(new_n561));
  XOR2_X1   g360(.A(KEYINPUT98), .B(KEYINPUT21), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G127gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n561), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n531), .B1(new_n567), .B2(KEYINPUT21), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G155gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  NOR4_X1   g380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(KEYINPUT100), .B(new_n577), .C1(new_n580), .C2(new_n581), .ZN(new_n583));
  INV_X1    g382(.A(G99gat), .ZN(new_n584));
  INV_X1    g383(.A(G106gat), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT8), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n583), .B(new_n586), .C1(G85gat), .C2(G92gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT101), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n589), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n593), .A2(new_n518), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n520), .B2(new_n593), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT99), .Z(new_n600));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT102), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(KEYINPUT102), .A3(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n576), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n588), .A2(KEYINPUT103), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(new_n590), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n590), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n560), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n567), .A2(new_n593), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n614), .A2(KEYINPUT10), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n609), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n618), .B2(new_n619), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT104), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n624), .B2(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n607), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n377), .A2(KEYINPUT105), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n377), .A2(KEYINPUT105), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n555), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  INV_X1    g437(.A(new_n460), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n555), .A2(new_n639), .A3(new_n632), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n640), .A2(G8gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT16), .B(G8gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT42), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(KEYINPUT42), .B2(new_n643), .ZN(G1325gat));
  NAND2_X1  g444(.A1(new_n555), .A2(new_n632), .ZN(new_n646));
  OAI21_X1  g445(.A(G15gat), .B1(new_n646), .B2(new_n476), .ZN(new_n647));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n555), .A2(new_n648), .A3(new_n470), .A4(new_n632), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(G1326gat));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n646), .B2(new_n488), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n555), .A2(KEYINPUT106), .A3(new_n416), .A4(new_n632), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  XOR2_X1   g455(.A(new_n576), .B(KEYINPUT108), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n547), .A2(new_n549), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n630), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT109), .ZN(new_n660));
  INV_X1    g459(.A(new_n606), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n504), .B2(new_n505), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n466), .A2(new_n503), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT110), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT110), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n466), .A2(new_n666), .A3(new_n503), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n606), .A2(KEYINPUT44), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n660), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G29gat), .B1(new_n671), .B2(new_n635), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n631), .A2(new_n576), .A3(new_n606), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n555), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n635), .A2(G29gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n673), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n675), .A2(new_n673), .A3(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n678), .A3(new_n679), .ZN(G1328gat));
  OAI21_X1  g479(.A(G36gat), .B1(new_n671), .B2(new_n460), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n460), .A2(G36gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT46), .B1(new_n675), .B2(new_n683), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n675), .A2(KEYINPUT46), .A3(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(G1329gat));
  AOI211_X1 g485(.A(new_n476), .B(new_n660), .C1(new_n663), .C2(new_n669), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT111), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n555), .A2(new_n688), .A3(new_n470), .A4(new_n674), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n687), .B2(new_n688), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OAI221_X1 g492(.A(new_n690), .B1(KEYINPUT111), .B2(KEYINPUT47), .C1(new_n687), .C2(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1330gat));
  AOI21_X1  g494(.A(new_n413), .B1(new_n670), .B2(new_n416), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n675), .A2(G50gat), .A3(new_n488), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1331gat));
  AND2_X1   g500(.A1(new_n665), .A2(new_n667), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n607), .A2(new_n658), .A3(new_n630), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n636), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n460), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT112), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n707), .A2(KEYINPUT113), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT113), .B1(new_n707), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n704), .A2(new_n715), .A3(new_n470), .ZN(new_n716));
  OAI21_X1  g515(.A(G71gat), .B1(new_n707), .B2(new_n476), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n416), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n576), .A2(new_n658), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n631), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n663), .B2(new_n669), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n635), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n606), .B1(new_n466), .B2(new_n503), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT114), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n722), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(KEYINPUT114), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n728), .A2(KEYINPUT114), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n722), .A4(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n636), .A2(new_n631), .A3(new_n580), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n726), .B1(new_n736), .B2(new_n737), .ZN(G1336gat));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n732), .A2(new_n739), .A3(new_n734), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT115), .B(new_n727), .C1(new_n730), .C2(new_n731), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n630), .A2(new_n460), .A3(G92gat), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n581), .B1(new_n724), .B2(new_n639), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT52), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n744), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT52), .B1(new_n735), .B2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n725), .B2(new_n476), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n631), .A2(new_n584), .A3(new_n470), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n736), .B2(new_n751), .ZN(G1338gat));
  NOR3_X1   g551(.A1(new_n630), .A2(G106gat), .A3(new_n488), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n740), .A2(new_n741), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n585), .B1(new_n724), .B2(new_n416), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT53), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n755), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT53), .B1(new_n735), .B2(new_n753), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1339gat));
  NAND3_X1  g559(.A1(new_n615), .A2(new_n609), .A3(new_n616), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n618), .A2(KEYINPUT54), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n622), .B1(new_n617), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT55), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT116), .Z(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(KEYINPUT55), .A3(new_n764), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n623), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n658), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n533), .A2(new_n534), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n537), .A2(new_n538), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n545), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT117), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n627), .A2(new_n773), .A3(new_n549), .A4(new_n629), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n661), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n766), .A2(new_n768), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n549), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n606), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n657), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n632), .A2(new_n547), .A3(new_n549), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n635), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n456), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n639), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(G113gat), .B1(new_n785), .B2(new_n658), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n416), .B1(new_n779), .B2(new_n780), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n639), .A2(new_n635), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n787), .A2(new_n470), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n554), .A2(new_n306), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(G1340gat));
  AOI21_X1  g590(.A(G120gat), .B1(new_n785), .B2(new_n631), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n630), .A2(new_n304), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n789), .B2(new_n793), .ZN(G1341gat));
  INV_X1    g593(.A(new_n789), .ZN(new_n795));
  OAI21_X1  g594(.A(G127gat), .B1(new_n795), .B2(new_n657), .ZN(new_n796));
  INV_X1    g595(.A(G127gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n785), .A2(new_n797), .A3(new_n576), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1342gat));
  OAI21_X1  g598(.A(G134gat), .B1(new_n795), .B2(new_n606), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n784), .A2(G134gat), .A3(new_n606), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n802), .A2(KEYINPUT118), .A3(new_n801), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT118), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  OAI221_X1 g603(.A(new_n800), .B1(new_n801), .B2(new_n802), .C1(new_n803), .C2(new_n804), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n476), .A2(new_n788), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n488), .B1(new_n779), .B2(new_n780), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n576), .ZN(new_n810));
  INV_X1    g609(.A(new_n778), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  INV_X1    g611(.A(new_n765), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n768), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n551), .B2(new_n552), .ZN(new_n815));
  INV_X1    g614(.A(new_n774), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n552), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n768), .B(new_n813), .C1(new_n818), .C2(new_n550), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(KEYINPUT119), .A3(new_n774), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n661), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n811), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT120), .B(new_n661), .C1(new_n817), .C2(new_n820), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n810), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n488), .B1(new_n825), .B2(new_n780), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n553), .B(new_n809), .C1(new_n826), .C2(new_n808), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G141gat), .ZN(new_n828));
  XOR2_X1   g627(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n829));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n781), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n781), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n476), .A2(new_n416), .A3(new_n460), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n553), .A2(new_n294), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT122), .Z(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n829), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n658), .B(new_n809), .C1(new_n826), .C2(new_n808), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n840), .A2(G141gat), .B1(new_n834), .B2(new_n837), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n292), .A2(KEYINPUT59), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n809), .B1(new_n826), .B2(new_n808), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n630), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n810), .B1(new_n821), .B2(new_n778), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n632), .A2(new_n554), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT57), .B(new_n488), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n779), .A2(new_n780), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n808), .B1(new_n850), .B2(new_n416), .ZN(new_n851));
  NOR4_X1   g650(.A1(new_n849), .A2(new_n630), .A3(new_n851), .A4(new_n806), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT59), .B1(new_n852), .B2(new_n292), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n834), .A2(new_n292), .A3(new_n631), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1345gat));
  OAI21_X1  g655(.A(G155gat), .B1(new_n845), .B2(new_n657), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n834), .A2(new_n298), .A3(new_n576), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1346gat));
  NAND2_X1  g658(.A1(new_n661), .A2(G162gat), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G162gat), .B1(new_n834), .B2(new_n661), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(G1347gat));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865));
  INV_X1    g664(.A(new_n787), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n636), .A2(new_n460), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n470), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n787), .A2(KEYINPUT125), .A3(new_n470), .A4(new_n867), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G169gat), .B1(new_n871), .B2(new_n554), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n782), .A2(new_n460), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT124), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n850), .A2(new_n635), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(KEYINPUT124), .B2(new_n873), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n227), .A3(new_n658), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n877), .ZN(G1348gat));
  OAI21_X1  g677(.A(G176gat), .B1(new_n871), .B2(new_n630), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n213), .A3(new_n631), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1349gat));
  OAI21_X1  g680(.A(G183gat), .B1(new_n871), .B2(new_n657), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n876), .A2(new_n238), .A3(new_n240), .A4(new_n576), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT60), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n882), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n876), .A2(new_n217), .A3(new_n661), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n661), .A3(new_n870), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(G190gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n217), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n891), .A2(new_n894), .B1(new_n890), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n893), .B2(new_n895), .ZN(G1351gat));
  INV_X1    g695(.A(new_n849), .ZN(new_n897));
  INV_X1    g696(.A(new_n851), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n476), .A2(new_n867), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n554), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n807), .A2(new_n900), .ZN(new_n904));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904), .B2(new_n658), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n905), .ZN(G1352gat));
  XOR2_X1   g705(.A(KEYINPUT127), .B(G204gat), .Z(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n631), .A3(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT62), .Z(new_n909));
  NOR2_X1   g708(.A1(new_n901), .A2(new_n630), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n907), .ZN(G1353gat));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n204), .A3(new_n576), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n576), .A3(new_n898), .A4(new_n900), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT63), .B1(new_n913), .B2(G211gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n901), .B2(new_n606), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n904), .A2(new_n205), .A3(new_n661), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1355gat));
endmodule


