//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G224), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT7), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(G128), .B(new_n194), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n200), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT0), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(new_n201), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n207), .A3(new_n201), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(new_n200), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n208), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n214), .A2(new_n215), .A3(new_n204), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n192), .B1(new_n206), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n208), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n212), .A2(new_n213), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n208), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n205), .B(new_n191), .C1(new_n220), .C2(new_n204), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G116), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT5), .ZN(new_n230));
  OAI21_X1  g044(.A(G113), .B1(new_n224), .B2(KEYINPUT5), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT88), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n225), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT5), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n236), .B(new_n237), .C1(new_n227), .C2(new_n235), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n229), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n241), .A2(KEYINPUT83), .A3(G107), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n241), .A2(KEYINPUT82), .A3(G107), .ZN(new_n245));
  INV_X1    g059(.A(G107), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G104), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G101), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n246), .A3(G104), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n244), .A2(new_n248), .A3(new_n249), .A4(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n241), .A2(G107), .ZN(new_n254));
  OAI21_X1  g068(.A(G101), .B1(new_n254), .B2(new_n247), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n239), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n230), .A2(new_n231), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n253), .B(new_n255), .C1(new_n229), .C2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT8), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n222), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n253), .A2(new_n255), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n239), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n248), .A2(new_n252), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT3), .B1(new_n251), .B2(KEYINPUT82), .ZN(new_n269));
  OAI21_X1  g083(.A(G101), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n270), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n272), .B(G101), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n227), .B(new_n228), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n267), .B(new_n260), .C1(new_n271), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n270), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n274), .A3(new_n273), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n280), .A2(KEYINPUT89), .A3(new_n267), .A4(new_n260), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n265), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n260), .B1(new_n280), .B2(new_n267), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT6), .ZN(new_n285));
  INV_X1    g099(.A(new_n284), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n273), .A2(new_n274), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n287), .A2(new_n279), .B1(new_n266), .B2(new_n239), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT89), .B1(new_n288), .B2(new_n260), .ZN(new_n289));
  INV_X1    g103(.A(new_n281), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n285), .B1(new_n291), .B2(KEYINPUT6), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n205), .B1(new_n220), .B2(new_n204), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n190), .B(KEYINPUT90), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n283), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT92), .ZN(new_n298));
  INV_X1    g112(.A(new_n285), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n284), .B1(new_n278), .B2(new_n281), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n295), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n283), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT93), .Z(new_n307));
  NAND3_X1  g121(.A1(new_n298), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n306), .A3(new_n283), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n188), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(KEYINPUT79), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(KEYINPUT79), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n196), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  OR3_X1    g130(.A1(new_n315), .A2(new_n204), .A3(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(G146), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT69), .A2(G237), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT69), .A2(G237), .ZN(new_n321));
  OAI211_X1 g135(.A(G214), .B(new_n189), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n193), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT69), .B(G237), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(G143), .A3(G214), .A4(new_n189), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT18), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n319), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(G131), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n327), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n316), .A2(KEYINPUT16), .A3(new_n317), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n204), .B2(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G146), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n196), .A3(new_n336), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n326), .B2(G131), .ZN(new_n342));
  AOI211_X1 g156(.A(KEYINPUT94), .B(new_n328), .C1(new_n323), .C2(new_n325), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n340), .B1(new_n344), .B2(KEYINPUT17), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT17), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n323), .A2(new_n325), .A3(new_n328), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n346), .B(new_n347), .C1(new_n342), .C2(new_n343), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n333), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G113), .B(G122), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(new_n241), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n331), .A2(KEYINPUT94), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n326), .A2(new_n341), .A3(G131), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT17), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n338), .A2(new_n339), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n348), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n330), .A2(new_n332), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n351), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT95), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT95), .A4(new_n351), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G475), .B1(new_n363), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n347), .B1(new_n342), .B2(new_n343), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT19), .B1(new_n312), .B2(new_n313), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n316), .A2(new_n317), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(KEYINPUT19), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n366), .B(new_n338), .C1(G146), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n351), .B1(new_n370), .B2(new_n358), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT95), .B1(new_n349), .B2(new_n351), .ZN(new_n373));
  INV_X1    g187(.A(new_n362), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(G475), .A2(G902), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n365), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n371), .B1(new_n361), .B2(new_n362), .ZN(new_n378));
  INV_X1    g192(.A(new_n376), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n378), .A2(KEYINPUT20), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n364), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(G234), .A2(G237), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n382), .A2(G952), .A3(new_n189), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n382), .A2(G902), .A3(G953), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT21), .B(G898), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G122), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT96), .B1(new_n387), .B2(G116), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n225), .A3(G122), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n225), .A2(G122), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(G107), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n193), .A2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n201), .A2(G143), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G134), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n391), .A2(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n388), .A2(new_n390), .A3(new_n400), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n394), .B(new_n399), .C1(new_n403), .C2(new_n246), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT13), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n395), .A2(KEYINPUT97), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(new_n396), .C1(new_n405), .C2(new_n395), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT97), .B1(new_n395), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g222(.A(G134), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n398), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n391), .A2(new_n392), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n246), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n409), .B(new_n410), .C1(new_n412), .C2(new_n393), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n415), .A2(new_n416), .A3(G953), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n404), .A2(new_n413), .A3(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G902), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n423), .B(new_n425), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n381), .A2(new_n386), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n189), .A2(G227), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND3_X1  g247(.A1(new_n279), .A2(new_n220), .A3(new_n273), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT68), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n198), .A2(new_n435), .A3(new_n202), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n198), .B2(new_n202), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT10), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n266), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n398), .A2(G137), .ZN(new_n441));
  AND2_X1   g255(.A1(KEYINPUT66), .A2(G137), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT66), .A2(G137), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n398), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n398), .B2(G137), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(KEYINPUT65), .B(new_n445), .C1(new_n398), .C2(G137), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n452), .A3(new_n328), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n198), .A2(new_n202), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n253), .A3(new_n255), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n434), .A2(new_n440), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n273), .A2(new_n220), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n464), .A2(new_n279), .B1(new_n439), .B2(new_n266), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n457), .A4(new_n461), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n456), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n433), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n473));
  INV_X1    g287(.A(new_n459), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n458), .B1(new_n253), .B2(new_n255), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n456), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n256), .A2(new_n203), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n459), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT12), .A4(new_n456), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT86), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n483), .A2(new_n484), .B1(new_n463), .B2(new_n467), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n473), .B1(new_n485), .B2(new_n433), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n482), .A3(new_n478), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n468), .A2(new_n487), .A3(new_n473), .A4(new_n433), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n472), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n422), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n468), .A2(new_n470), .A3(new_n433), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n485), .B2(new_n433), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n491), .B1(new_n494), .B2(new_n422), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n430), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n310), .A2(new_n428), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n223), .B2(G128), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n500), .A2(KEYINPUT23), .B1(new_n223), .B2(G128), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT23), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n499), .B(new_n502), .C1(new_n223), .C2(G128), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G110), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT76), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  XNOR2_X1  g322(.A(G119), .B(G128), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n340), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT78), .B(G110), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n504), .A2(new_n512), .B1(new_n509), .B2(new_n508), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n338), .A2(new_n513), .A3(new_n314), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT22), .B(G137), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n515), .B(new_n516), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n511), .B2(new_n514), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n422), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT25), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n422), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n416), .B1(G234), .B2(new_n422), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT81), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT80), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n520), .B2(new_n521), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n511), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n517), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT80), .A3(new_n519), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n526), .A2(G902), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  AOI211_X1 g351(.A(KEYINPUT81), .B(new_n537), .C1(new_n530), .C2(new_n533), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n527), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G472), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n324), .A2(G210), .A3(new_n189), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n542), .B(new_n543), .Z(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n447), .A2(new_n452), .A3(new_n328), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n328), .B1(new_n447), .B2(new_n452), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n220), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n444), .A2(G134), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n398), .A2(G137), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n198), .A2(new_n435), .A3(new_n202), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n551), .A2(new_n554), .A3(new_n455), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT71), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n550), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n274), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT28), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n455), .A2(new_n554), .A3(new_n458), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT67), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n554), .A2(new_n455), .A3(new_n458), .A4(KEYINPUT67), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n550), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n274), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n550), .A2(new_n556), .A3(new_n562), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n564), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n547), .B1(new_n563), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n571), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT30), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n567), .A2(new_n576), .A3(new_n550), .A4(new_n568), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n578), .B2(new_n274), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n546), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n579), .B2(new_n546), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n541), .B(new_n422), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT32), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n546), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT31), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n581), .A3(new_n573), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n541), .A4(new_n422), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n550), .A2(new_n559), .A3(new_n556), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n559), .B1(new_n550), .B2(new_n556), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n562), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n564), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n557), .A2(new_n274), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n571), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT28), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n546), .A2(KEYINPUT29), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n422), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n456), .A2(new_n220), .B1(new_n565), .B2(new_n566), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n562), .B1(new_n602), .B2(new_n568), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT28), .B1(new_n603), .B2(new_n574), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n595), .A3(new_n546), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT72), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n604), .A2(new_n595), .A3(KEYINPUT72), .A4(new_n546), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n578), .A2(new_n274), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n571), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT29), .B1(new_n610), .B2(new_n547), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n601), .B1(new_n612), .B2(KEYINPUT73), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n607), .A2(new_n611), .A3(new_n614), .A4(new_n608), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n541), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT74), .B1(new_n591), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(KEYINPUT73), .ZN(new_n618));
  INV_X1    g432(.A(new_n601), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT74), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n585), .A2(new_n590), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n498), .A2(new_n540), .A3(new_n617), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT98), .B(G101), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G3));
  INV_X1    g441(.A(new_n584), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n541), .B1(new_n588), .B2(new_n422), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n539), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n497), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  INV_X1    g446(.A(new_n306), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n297), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n188), .B1(new_n634), .B2(new_n309), .ZN(new_n635));
  INV_X1    g449(.A(new_n386), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n420), .A2(KEYINPUT101), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n404), .A2(new_n639), .A3(new_n413), .A4(new_n417), .ZN(new_n640));
  AND4_X1   g454(.A1(KEYINPUT33), .A2(new_n638), .A3(new_n419), .A4(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT33), .B1(new_n419), .B2(new_n420), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n424), .A2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT102), .B(G478), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n423), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n381), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n637), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT103), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND3_X1  g470(.A1(new_n375), .A2(new_n365), .A3(new_n376), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT20), .B1(new_n378), .B2(new_n379), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n427), .A3(new_n364), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n637), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n632), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n518), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n531), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n535), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n527), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n669), .A2(new_n628), .A3(new_n629), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n310), .A2(new_n670), .A3(new_n497), .A4(new_n428), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  AND3_X1   g487(.A1(new_n303), .A2(new_n306), .A3(new_n283), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n306), .B1(new_n303), .B2(new_n283), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n668), .B(new_n187), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n384), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n383), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n676), .A2(new_n660), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n617), .A2(new_n624), .A3(new_n497), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XOR2_X1   g498(.A(new_n680), .B(KEYINPUT39), .Z(new_n685));
  AOI211_X1 g499(.A(new_n430), .B(new_n685), .C1(new_n492), .C2(new_n496), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n308), .A2(new_n309), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n691));
  XOR2_X1   g505(.A(new_n690), .B(new_n691), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n597), .A2(new_n547), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT105), .Z(new_n694));
  INV_X1    g508(.A(new_n586), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n422), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n623), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n426), .B1(new_n659), .B2(new_n364), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n187), .A2(new_n698), .A3(new_n669), .A4(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n688), .A2(new_n689), .A3(new_n692), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  NAND3_X1  g516(.A1(new_n381), .A2(new_n650), .A3(new_n680), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n676), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n617), .A2(new_n624), .A3(new_n497), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NOR3_X1   g520(.A1(new_n591), .A2(new_n616), .A3(KEYINPUT74), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n468), .A2(new_n433), .A3(new_n487), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT87), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n471), .B1(new_n711), .B2(new_n488), .ZN(new_n712));
  OAI21_X1  g526(.A(G469), .B1(new_n712), .B2(G902), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n492), .A2(new_n713), .A3(new_n429), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n492), .A2(new_n713), .A3(KEYINPUT106), .A4(new_n429), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n709), .A2(new_n540), .A3(new_n652), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n709), .A2(new_n540), .A3(new_n661), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AND3_X1   g537(.A1(new_n716), .A2(new_n635), .A3(new_n717), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n381), .A2(new_n669), .A3(new_n386), .A4(new_n427), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n709), .A2(new_n724), .A3(KEYINPUT107), .A4(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n617), .A2(new_n624), .A3(new_n725), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n716), .A2(new_n635), .A3(new_n717), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NAND2_X1  g546(.A1(new_n588), .A2(new_n422), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT108), .B(G472), .Z(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(G472), .A2(G902), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n595), .A2(new_n598), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n581), .B1(new_n738), .B2(new_n546), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n739), .B2(new_n583), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n736), .A2(new_n741), .A3(new_n539), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n635), .A2(new_n699), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n636), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n716), .A2(new_n717), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n387), .ZN(G24));
  OAI211_X1 g561(.A(new_n740), .B(new_n668), .C1(new_n734), .C2(new_n735), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n703), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n716), .A3(new_n635), .A4(new_n717), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  INV_X1    g565(.A(new_n703), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n712), .A2(G469), .A3(G902), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT109), .B1(new_n753), .B2(new_n495), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n492), .A2(new_n496), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n308), .A2(new_n187), .A3(new_n309), .A4(new_n429), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n709), .A2(new_n540), .A3(new_n752), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n621), .A2(new_n623), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n381), .A2(new_n650), .A3(KEYINPUT42), .A4(new_n680), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n540), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n307), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n297), .B2(KEYINPUT92), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n188), .B(new_n674), .C1(new_n768), .C2(new_n305), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n429), .A3(new_n754), .A4(new_n756), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n762), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n620), .A2(G472), .B1(new_n585), .B2(new_n590), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n772), .A2(new_n539), .A3(new_n764), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n759), .A2(new_n773), .A3(KEYINPUT110), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n760), .A2(new_n761), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT111), .B(G131), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G33));
  NOR2_X1   g591(.A1(new_n660), .A2(new_n681), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n709), .A2(new_n540), .A3(new_n778), .A4(new_n759), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  XNOR2_X1  g594(.A(new_n494), .B(KEYINPUT45), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(G469), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n491), .A2(new_n422), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n753), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(KEYINPUT46), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n429), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n685), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n308), .A2(new_n187), .A3(new_n309), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n373), .A2(new_n374), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n422), .B1(new_n790), .B2(new_n352), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n657), .A2(new_n658), .B1(new_n791), .B2(G475), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n650), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT43), .Z(new_n794));
  OAI21_X1  g608(.A(new_n668), .B1(new_n628), .B2(new_n629), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n789), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n788), .B(new_n801), .C1(new_n800), .C2(new_n799), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NOR4_X1   g617(.A1(new_n709), .A2(new_n540), .A3(new_n703), .A4(new_n789), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n786), .A2(KEYINPUT47), .A3(new_n429), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n786), .B2(new_n429), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  INV_X1    g623(.A(new_n742), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n794), .A2(new_n383), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n794), .A2(new_n813), .A3(new_n383), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n810), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n769), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n805), .A2(new_n806), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n492), .A2(new_n713), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n429), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n817), .B2(KEYINPUT117), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n812), .A2(new_n814), .ZN(new_n823));
  INV_X1    g637(.A(new_n748), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n745), .A2(new_n789), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n698), .A2(new_n539), .A3(new_n679), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n792), .A2(new_n647), .A3(new_n649), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n692), .A2(new_n187), .A3(new_n745), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT50), .B1(new_n815), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n809), .B1(new_n822), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n763), .A2(new_n540), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n823), .A2(new_n840), .A3(new_n825), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT120), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n844), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n842), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT48), .ZN(new_n849));
  OAI211_X1 g663(.A(G952), .B(new_n189), .C1(new_n828), .C2(new_n651), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n815), .B2(new_n724), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT48), .ZN(new_n852));
  OAI211_X1 g666(.A(KEYINPUT120), .B(new_n852), .C1(new_n843), .C2(new_n844), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n838), .A2(new_n849), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n668), .A2(new_n430), .A3(new_n681), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n855), .A2(new_n635), .A3(new_n699), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n698), .A3(new_n754), .A4(new_n756), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n683), .A2(new_n705), .A3(new_n750), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT52), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n683), .A2(new_n705), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT115), .A3(new_n750), .A4(new_n857), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n858), .A2(new_n859), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n617), .A2(new_n540), .A3(new_n624), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n745), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n746), .B1(new_n870), .B2(new_n652), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n731), .A3(new_n872), .A4(new_n722), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n386), .B1(new_n651), .B2(new_n660), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n310), .A3(new_n497), .A4(new_n630), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n875), .A2(new_n671), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n876), .A2(new_n625), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n726), .A2(new_n730), .ZN(new_n879));
  INV_X1    g693(.A(new_n746), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n719), .A2(new_n722), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT114), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n792), .A2(new_n426), .A3(new_n668), .A4(new_n680), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n789), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n617), .A2(new_n884), .A3(new_n624), .A4(new_n497), .ZN(new_n885));
  INV_X1    g699(.A(new_n758), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n749), .A2(new_n886), .A3(new_n754), .A4(new_n756), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n779), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n775), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n868), .A2(new_n878), .A3(new_n882), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT53), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n858), .A2(new_n865), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n867), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n882), .A2(new_n889), .A3(new_n873), .A4(new_n877), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n897), .A3(KEYINPUT54), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n876), .A2(new_n625), .A3(KEYINPUT53), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n871), .A3(new_n731), .A4(new_n722), .ZN(new_n900));
  INV_X1    g714(.A(new_n778), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n869), .A2(new_n901), .A3(new_n770), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n885), .A2(new_n887), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n869), .A2(new_n770), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT42), .B1(new_n905), .B2(new_n752), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n771), .A2(new_n774), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n893), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n890), .B2(new_n894), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n836), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n831), .B1(new_n914), .B2(new_n834), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(KEYINPUT118), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n832), .B(KEYINPUT118), .C1(new_n835), .C2(new_n836), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n817), .B1(new_n429), .B2(new_n819), .ZN(new_n918));
  INV_X1    g732(.A(new_n816), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n809), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n854), .A2(new_n898), .A3(new_n913), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(G952), .B2(G953), .ZN(new_n923));
  INV_X1    g737(.A(new_n692), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT113), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n540), .A2(new_n187), .A3(new_n429), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n698), .A2(new_n928), .A3(new_n793), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n924), .A2(new_n926), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n923), .A2(new_n930), .ZN(G75));
  XNOR2_X1  g745(.A(new_n302), .B(new_n296), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n911), .A2(new_n422), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n633), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n189), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n911), .A2(new_n422), .A3(new_n767), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n933), .A2(new_n936), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n937), .A2(new_n942), .ZN(G51));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n862), .A2(new_n867), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n894), .B1(new_n945), .B2(new_n896), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n909), .A2(new_n893), .ZN(new_n947));
  AND4_X1   g761(.A1(new_n944), .A2(new_n946), .A3(new_n912), .A4(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n911), .B2(new_n912), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n913), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n783), .B(KEYINPUT57), .Z(new_n951));
  OAI21_X1  g765(.A(new_n490), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n934), .A2(new_n782), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n938), .B1(new_n952), .B2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n378), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n378), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n938), .ZN(G60));
  INV_X1    g772(.A(new_n645), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  NOR3_X1   g775(.A1(new_n950), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n913), .B2(new_n898), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n939), .B1(new_n963), .B2(new_n645), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT122), .Z(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT60), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n946), .B2(new_n947), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n939), .B1(new_n970), .B2(new_n534), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n666), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n977));
  INV_X1    g791(.A(new_n974), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n976), .B(new_n977), .C1(new_n978), .C2(new_n971), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n975), .A2(new_n979), .ZN(G66));
  NAND2_X1  g794(.A1(new_n878), .A2(new_n882), .ZN(new_n981));
  NAND2_X1  g795(.A1(G224), .A2(G953), .ZN(new_n982));
  OAI22_X1  g796(.A1(new_n981), .A2(G953), .B1(new_n385), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n292), .B1(G898), .B2(new_n189), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT124), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  XNOR2_X1  g800(.A(new_n578), .B(KEYINPUT125), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(new_n369), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n802), .A2(new_n807), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n789), .B1(new_n651), .B2(new_n660), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n709), .A2(new_n540), .A3(new_n686), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n863), .A2(new_n750), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n701), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n989), .B1(new_n997), .B2(G953), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n999));
  INV_X1    g813(.A(new_n775), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n840), .A2(new_n743), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n902), .B1(new_n788), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n990), .A2(new_n1000), .A3(new_n994), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n998), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G72));
  NAND3_X1  g821(.A1(new_n997), .A2(new_n882), .A3(new_n878), .ZN(new_n1008));
  XNOR2_X1  g822(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n541), .A2(new_n422), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n610), .B(KEYINPUT127), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n546), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n610), .A2(new_n547), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n586), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n891), .A2(new_n897), .A3(new_n1011), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1011), .B1(new_n1003), .B2(new_n981), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1013), .A2(new_n546), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n938), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1014), .A2(new_n1017), .A3(new_n1020), .ZN(G57));
endmodule


