//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(G952), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AOI211_X1 g008(.A(new_n193), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT21), .B(G898), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT80), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(KEYINPUT80), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n199), .A2(new_n202), .A3(KEYINPUT80), .A4(G104), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n207), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT68), .A2(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT68), .A2(G116), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G119), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n216), .B(new_n221), .C1(new_n222), .C2(G119), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n222), .A2(G119), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n217), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n216), .B1(new_n222), .B2(G119), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n224), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n213), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n206), .A2(G107), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n208), .A2(new_n207), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n219), .A2(G113), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(new_n215), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT68), .A2(G116), .ZN(new_n244));
  INV_X1    g058(.A(G119), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n241), .B(new_n242), .C1(new_n246), .C2(new_n225), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(G101), .C1(new_n234), .C2(new_n235), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n237), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G122), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n229), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n228), .A2(new_n212), .A3(new_n223), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(KEYINPUT8), .ZN(new_n255));
  INV_X1    g069(.A(new_n223), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n216), .B(KEYINPUT5), .C1(new_n222), .C2(G119), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n226), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n254), .B(new_n255), .C1(new_n258), .C2(new_n212), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT87), .ZN(new_n260));
  INV_X1    g074(.A(G224), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n194), .A2(KEYINPUT87), .A3(G224), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(KEYINPUT65), .A3(G146), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(G143), .B2(new_n271), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n265), .A2(KEYINPUT64), .A3(G146), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n268), .B(new_n269), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(G143), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(new_n266), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n274), .A2(new_n277), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G125), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n265), .A2(KEYINPUT65), .A3(G146), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT65), .B1(new_n265), .B2(G146), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT64), .B1(new_n265), .B2(G146), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n270), .A2(new_n271), .A3(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G128), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n285), .A2(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n278), .A2(new_n266), .A3(new_n296), .A4(G128), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n295), .A2(G125), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n264), .B1(new_n282), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n274), .A2(new_n277), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n279), .A2(new_n275), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n293), .A2(new_n294), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n274), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n281), .ZN(new_n307));
  INV_X1    g121(.A(new_n264), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n253), .A2(new_n259), .A3(new_n300), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n193), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT88), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n229), .A2(new_n251), .ZN(new_n313));
  INV_X1    g127(.A(new_n252), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT6), .A3(new_n253), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n307), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n262), .A2(new_n263), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT86), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT6), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n313), .A2(new_n321), .A3(new_n314), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G210), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n310), .A2(new_n325), .A3(new_n193), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n312), .A2(new_n323), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n324), .B(KEYINPUT90), .Z(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n312), .A2(new_n323), .A3(new_n326), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n312), .A2(new_n323), .A3(KEYINPUT89), .A4(new_n326), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G214), .B1(G237), .B2(G902), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT92), .B(G104), .Z(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT74), .A2(G140), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT74), .A2(G140), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n341), .B(G125), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OR2_X1    g158(.A1(KEYINPUT74), .A2(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT74), .A2(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n281), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n281), .A2(G140), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT75), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n344), .B(KEYINPUT19), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G125), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(new_n348), .ZN(new_n353));
  OR2_X1    g167(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n271), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n344), .B(KEYINPUT16), .C1(new_n347), .C2(new_n349), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G146), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n190), .A2(new_n194), .A3(G214), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(new_n265), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G131), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n364), .B(G143), .ZN(new_n367));
  INV_X1    g181(.A(G131), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT18), .A2(G131), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n365), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n271), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n344), .B1(new_n347), .B2(new_n349), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(new_n271), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n340), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT17), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n359), .A2(new_n271), .A3(new_n361), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n365), .A2(KEYINPUT17), .A3(G131), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n381), .A2(new_n363), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n377), .A3(new_n340), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n385), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT20), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n340), .B1(new_n384), .B2(new_n377), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n193), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n214), .A2(G122), .A3(new_n215), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n222), .B2(G122), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n214), .A2(new_n399), .A3(G122), .A4(new_n215), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n402), .A2(KEYINPUT94), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(G107), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n398), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n222), .A2(G122), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n408), .A2(G107), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n290), .A2(new_n292), .A3(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n265), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G134), .ZN(new_n414));
  INV_X1    g228(.A(G134), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n410), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(KEYINPUT93), .A3(new_n416), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT95), .A4(G107), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n407), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT13), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n411), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n413), .A3(G134), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n423), .A2(new_n415), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n408), .A2(new_n409), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n202), .ZN(new_n428));
  OAI221_X1 g242(.A(new_n425), .B1(new_n413), .B2(new_n426), .C1(new_n428), .C2(new_n410), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  INV_X1    g244(.A(G217), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(G953), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n422), .B2(new_n429), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n193), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT96), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT15), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n422), .A2(new_n429), .ZN(new_n440));
  INV_X1    g254(.A(new_n432), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n433), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n193), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n442), .B2(new_n433), .ZN(new_n448));
  INV_X1    g262(.A(new_n439), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n437), .A2(new_n445), .A3(new_n447), .A4(new_n439), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n397), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND4_X1   g267(.A1(new_n198), .A2(new_n336), .A3(new_n337), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT32), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT11), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n415), .B2(G137), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT11), .A3(G134), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n415), .A2(G137), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n368), .A4(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n415), .A2(G137), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n458), .A2(G134), .ZN(new_n463));
  OAI21_X1  g277(.A(G131), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n295), .B2(new_n298), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n301), .A3(new_n302), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n466), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n248), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n247), .A2(new_n475), .A3(new_n223), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n247), .B2(new_n223), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n466), .A2(new_n470), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT70), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n248), .A2(KEYINPUT69), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n247), .A2(new_n475), .A3(new_n223), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n274), .A2(new_n305), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n297), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n485), .A2(new_n465), .B1(new_n280), .B2(new_n469), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n190), .A2(new_n194), .A3(G210), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT27), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT26), .B(G101), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n474), .A2(new_n480), .A3(new_n488), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT31), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n479), .A2(new_n248), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n495), .A3(new_n488), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT28), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT28), .B1(new_n483), .B2(new_n486), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n492), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(G472), .A2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n455), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n493), .B(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n496), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT71), .B1(new_n496), .B2(KEYINPUT28), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n511), .A2(new_n512), .A3(new_n501), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n510), .B1(new_n513), .B2(new_n492), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(KEYINPUT32), .A3(new_n506), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n478), .A2(new_n479), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n480), .A2(new_n488), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT28), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n501), .A2(new_n520), .A3(new_n504), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n193), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n501), .A2(new_n504), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n511), .A2(new_n512), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n474), .A2(new_n480), .A3(new_n488), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT29), .B1(new_n528), .B2(new_n504), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n524), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n531), .B2(G472), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n499), .A2(new_n500), .A3(new_n525), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n523), .B1(new_n533), .B2(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(G472), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n534), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n508), .B(new_n515), .C1(new_n532), .C2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT22), .B(G137), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n538), .B(new_n539), .Z(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n363), .A2(new_n382), .ZN(new_n542));
  AND2_X1   g356(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n543));
  NOR2_X1   g357(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n544));
  OAI22_X1  g358(.A1(new_n543), .A2(new_n544), .B1(new_n245), .B2(G128), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n289), .A2(G119), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n290), .A2(new_n292), .A3(G119), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT23), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n545), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G110), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT66), .B(G128), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n546), .B1(new_n552), .B2(G119), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT24), .B(G110), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n542), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT76), .B1(new_n553), .B2(new_n555), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(KEYINPUT23), .A3(G119), .ZN(new_n561));
  INV_X1    g375(.A(G110), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n545), .A3(new_n562), .A4(new_n547), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n548), .A2(new_n547), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n554), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n363), .A2(new_n567), .A3(new_n374), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n541), .B1(new_n559), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT77), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n363), .A2(new_n567), .A3(new_n374), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n557), .B1(new_n363), .B2(new_n382), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n559), .A2(KEYINPUT77), .A3(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n569), .B1(new_n575), .B2(new_n541), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n189), .B2(G217), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G217), .B1(new_n189), .B2(G902), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT78), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n576), .B2(G902), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n582), .B(KEYINPUT25), .C1(new_n576), .C2(G902), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n289), .B1(new_n278), .B2(KEYINPUT1), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n297), .B1(new_n279), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n590), .A2(new_n209), .A3(new_n211), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n213), .A2(new_n485), .A3(KEYINPUT10), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n237), .A2(new_n250), .A3(new_n280), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n469), .B(KEYINPUT81), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(G110), .B(G140), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT79), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n194), .A2(G227), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n598), .B(new_n599), .Z(new_n600));
  AND2_X1   g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n469), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n212), .A2(new_n306), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT82), .ZN(new_n606));
  INV_X1    g420(.A(new_n591), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT82), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n212), .A2(new_n306), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n610), .A2(KEYINPUT12), .A3(new_n469), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT12), .B1(new_n610), .B2(new_n469), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT83), .B(new_n596), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n600), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT12), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n212), .A2(new_n306), .A3(new_n608), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n608), .B1(new_n212), .B2(new_n306), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n617), .A2(new_n618), .A3(new_n591), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n602), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(KEYINPUT12), .A3(new_n469), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT83), .B1(new_n622), .B2(new_n596), .ZN(new_n623));
  OAI211_X1 g437(.A(G469), .B(new_n604), .C1(new_n615), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G469), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n193), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT84), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n611), .B2(new_n612), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n620), .A2(KEYINPUT84), .A3(new_n621), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n601), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n596), .B1(new_n603), .B2(new_n602), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n614), .ZN(new_n634));
  AOI211_X1 g448(.A(G469), .B(G902), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n588), .B1(new_n628), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n454), .A2(new_n537), .A3(new_n587), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n535), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n505), .A2(G902), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n641), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n514), .B2(new_n193), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n637), .A3(new_n587), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n437), .A2(new_n438), .A3(new_n445), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n438), .A2(G902), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n443), .A2(KEYINPUT33), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n442), .B2(new_n433), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n648), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n198), .A3(new_n397), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n655));
  INV_X1    g469(.A(new_n324), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n331), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n327), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n658), .B2(new_n337), .ZN(new_n659));
  INV_X1    g473(.A(new_n337), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT99), .B(new_n660), .C1(new_n657), .C2(new_n327), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n654), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n646), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT34), .B(G104), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n393), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT100), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n668), .A2(new_n669), .B1(G475), .B2(new_n395), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n198), .A3(new_n451), .A4(new_n452), .ZN(new_n671));
  OR3_X1    g485(.A1(new_n671), .A2(new_n661), .A3(new_n659), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n646), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT35), .B(G107), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n585), .A2(new_n586), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n575), .B(new_n677), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n578), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n454), .A2(new_n637), .A3(new_n645), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NOR3_X1   g497(.A1(new_n636), .A2(new_n661), .A3(new_n659), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n192), .B1(new_n195), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n670), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n451), .A2(new_n452), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n684), .A2(new_n537), .A3(new_n680), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n680), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n505), .A2(new_n455), .A3(new_n507), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT32), .B1(new_n514), .B2(new_n506), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n531), .A2(new_n516), .A3(G472), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT72), .B1(new_n534), .B2(new_n535), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n694), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(KEYINPUT101), .A3(new_n690), .A4(new_n684), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  NAND2_X1  g518(.A1(new_n336), .A2(KEYINPUT38), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n335), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n451), .A2(new_n397), .A3(new_n452), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n680), .A2(new_n660), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n518), .A2(new_n492), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n528), .A2(new_n492), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(KEYINPUT102), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n193), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT102), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n508), .A2(new_n515), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n708), .A2(new_n710), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n686), .B(KEYINPUT39), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n637), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT40), .Z(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n722), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  AND3_X1   g539(.A1(new_n653), .A2(new_n397), .A3(new_n687), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n684), .A2(new_n537), .A3(new_n680), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT104), .B(G146), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G48));
  INV_X1    g543(.A(new_n587), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n697), .B2(new_n700), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n632), .A2(new_n634), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n625), .B1(new_n732), .B2(new_n193), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n635), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT105), .B1(new_n734), .B2(new_n588), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  INV_X1    g550(.A(new_n588), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n733), .A2(new_n635), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n731), .A2(new_n662), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NOR3_X1   g556(.A1(new_n671), .A2(new_n661), .A3(new_n659), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n731), .A2(new_n743), .A3(new_n739), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  AND2_X1   g559(.A1(new_n632), .A2(new_n634), .ZN(new_n746));
  OAI21_X1  g560(.A(G469), .B1(new_n746), .B2(G902), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n732), .A2(new_n625), .A3(new_n193), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n588), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n661), .A3(new_n659), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n453), .A2(new_n198), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n537), .A3(new_n680), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  XOR2_X1   g567(.A(KEYINPUT106), .B(G472), .Z(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n505), .B2(G902), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n492), .B1(new_n519), .B2(new_n502), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n506), .B1(new_n494), .B2(new_n756), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n198), .A2(new_n755), .A3(new_n587), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n749), .A2(new_n736), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n659), .A2(new_n661), .A3(new_n709), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n734), .A2(KEYINPUT105), .A3(new_n588), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  AND4_X1   g577(.A1(new_n680), .A2(new_n726), .A3(new_n757), .A4(new_n755), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n750), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NAND2_X1  g580(.A1(new_n335), .A2(new_n337), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n636), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n537), .A2(new_n768), .A3(new_n587), .A4(new_n726), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n731), .A2(new_n726), .A3(new_n768), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  NAND4_X1  g592(.A1(new_n537), .A2(new_n768), .A3(new_n690), .A4(new_n587), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n731), .A2(new_n781), .A3(new_n690), .A4(new_n768), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  INV_X1    g598(.A(new_n397), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n653), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT43), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n397), .B1(new_n647), .B2(new_n652), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n680), .C1(new_n644), .C2(new_n642), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n767), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n795), .B(new_n796), .C1(new_n794), .C2(new_n792), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n604), .B1(new_n615), .B2(new_n623), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n625), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT45), .B(new_n604), .C1(new_n615), .C2(new_n623), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n626), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n748), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n805), .A2(KEYINPUT46), .A3(new_n627), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n588), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n719), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n797), .A2(new_n798), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n458), .ZN(G39));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT47), .B(new_n588), .C1(new_n804), .C2(new_n806), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n796), .A2(new_n730), .A3(new_n726), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n537), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  INV_X1    g633(.A(new_n764), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n689), .A2(new_n670), .A3(new_n687), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n537), .A2(new_n680), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n768), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n777), .A2(new_n783), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n740), .A2(new_n638), .A3(new_n681), .A4(new_n752), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n654), .A2(new_n335), .A3(new_n660), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n645), .A2(new_n827), .A3(new_n637), .A4(new_n587), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n537), .A2(new_n759), .A3(new_n587), .A4(new_n761), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n762), .B(new_n828), .C1(new_n829), .C2(new_n672), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n335), .A2(new_n197), .A3(new_n660), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n689), .A2(new_n397), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n831), .A2(KEYINPUT111), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT111), .B1(new_n831), .B2(new_n832), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n646), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n826), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n825), .A2(new_n836), .A3(KEYINPUT53), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n680), .A2(new_n686), .A3(new_n709), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n684), .A2(new_n839), .A3(new_n717), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n727), .A2(new_n765), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n703), .A2(new_n841), .A3(KEYINPUT52), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(new_n703), .B2(new_n841), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n703), .A2(new_n841), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n703), .A2(new_n841), .A3(KEYINPUT52), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n838), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  XNOR2_X1  g666(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n842), .A2(new_n843), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n825), .A2(new_n836), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n830), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n740), .A2(new_n681), .ZN(new_n861));
  INV_X1    g675(.A(new_n835), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n638), .A2(new_n752), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n777), .A2(new_n783), .A3(new_n824), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n848), .A2(new_n849), .ZN(new_n867));
  INV_X1    g681(.A(new_n853), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT112), .B1(new_n842), .B2(new_n843), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n848), .A2(new_n845), .A3(new_n849), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n855), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n869), .B1(new_n872), .B2(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n851), .A2(new_n856), .A3(KEYINPUT114), .A4(new_n852), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n734), .A2(KEYINPUT115), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n734), .A2(KEYINPUT115), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n737), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n813), .A2(new_n814), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n787), .A2(new_n790), .A3(new_n192), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n755), .A2(new_n757), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n587), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n767), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n747), .A2(new_n748), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n588), .A2(new_n192), .A3(new_n337), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n336), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n697), .A3(new_n587), .A4(new_n716), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n785), .A2(new_n647), .A3(new_n652), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n791), .A2(new_n888), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n882), .A2(new_n680), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n889), .A2(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT50), .ZN(new_n894));
  INV_X1    g708(.A(new_n749), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n705), .A3(new_n660), .A4(new_n707), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n883), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n896), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n882), .A2(new_n587), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(KEYINPUT50), .A3(new_n899), .A4(new_n881), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n893), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT51), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n885), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n731), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n891), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT48), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n899), .A2(new_n750), .A3(new_n881), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n653), .A2(new_n397), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n188), .C1(new_n912), .C2(new_n889), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n876), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n885), .A2(new_n901), .A3(new_n904), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n904), .B1(new_n885), .B2(new_n901), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n876), .B(new_n914), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n859), .A2(new_n874), .A3(new_n875), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT117), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n837), .B1(new_n870), .B2(new_n871), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT54), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n925), .A2(KEYINPUT114), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT117), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n859), .A4(new_n920), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n187), .A2(new_n194), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n922), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n587), .A2(new_n788), .A3(new_n337), .A4(new_n588), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT110), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n886), .B(KEYINPUT49), .ZN(new_n933));
  OR4_X1    g747(.A1(new_n708), .A2(new_n932), .A3(new_n717), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G75));
  OAI211_X1 g749(.A(G210), .B(G902), .C1(new_n923), .C2(new_n924), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n316), .A2(new_n322), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n320), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT55), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n194), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(G902), .B(new_n329), .C1(new_n923), .C2(new_n924), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n942), .B(new_n944), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT120), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n943), .B1(new_n938), .B2(new_n941), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n953), .B(new_n954), .C1(new_n950), .C2(new_n949), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(G51));
  OAI21_X1  g770(.A(KEYINPUT54), .B1(new_n923), .B2(new_n924), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n857), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n626), .B(KEYINPUT57), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n746), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n805), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n193), .B1(new_n851), .B2(new_n856), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n960), .A2(KEYINPUT121), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT121), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n958), .A2(new_n959), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n746), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n943), .B1(new_n963), .B2(new_n966), .ZN(G54));
  NAND3_X1  g781(.A1(new_n962), .A2(KEYINPUT58), .A3(G475), .ZN(new_n968));
  INV_X1    g782(.A(new_n386), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(new_n943), .ZN(G60));
  INV_X1    g786(.A(new_n958), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n649), .A2(new_n651), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT59), .Z(new_n977));
  OR2_X1    g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n944), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n926), .A2(new_n859), .ZN(new_n980));
  INV_X1    g794(.A(new_n977), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n982), .B2(new_n975), .ZN(G63));
  NAND2_X1  g797(.A1(new_n851), .A2(new_n856), .ZN(new_n984));
  XNOR2_X1  g798(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n431), .A2(new_n193), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n678), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n984), .A2(new_n987), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n944), .B(new_n988), .C1(new_n989), .C2(new_n577), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G66));
  INV_X1    g806(.A(new_n196), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n194), .B1(new_n993), .B2(G224), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n864), .B2(new_n194), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n939), .B1(G898), .B2(new_n194), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT124), .Z(new_n997));
  XNOR2_X1  g811(.A(new_n995), .B(new_n997), .ZN(G69));
  AOI21_X1  g812(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n810), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n808), .A2(new_n719), .A3(new_n731), .A4(new_n760), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n777), .A2(new_n783), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1001), .A2(new_n1002), .A3(new_n818), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n703), .A2(new_n727), .A3(new_n765), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1004), .A2(G953), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n472), .A2(new_n473), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n357), .B(KEYINPUT125), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n685), .B2(new_n194), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1009), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n724), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n796), .B1(new_n911), .B2(new_n832), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n907), .A2(new_n720), .A3(new_n1020), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n1021), .B(new_n810), .C1(new_n815), .C2(new_n817), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT62), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1017), .A2(new_n1023), .A3(new_n724), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1025), .A2(new_n194), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1000), .B(new_n1016), .C1(new_n1026), .C2(new_n1013), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1013), .B1(new_n1025), .B2(new_n194), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n999), .B1(new_n1028), .B2(new_n1015), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(G72));
  NAND4_X1  g844(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .A4(new_n836), .ZN(new_n1031));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  AOI21_X1  g847(.A(new_n712), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1004), .A2(new_n1009), .A3(new_n864), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1033), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1037), .A2(new_n492), .A3(new_n528), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n528), .A2(new_n504), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT127), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1036), .B1(new_n1040), .B2(new_n493), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n873), .A2(new_n1041), .ZN(new_n1042));
  NOR4_X1   g856(.A1(new_n1034), .A2(new_n1038), .A3(new_n943), .A4(new_n1042), .ZN(G57));
endmodule


