//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n203), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n214), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n204), .A2(new_n205), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n212), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n217), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G33), .A3(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n231), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G226), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n258), .A2(G274), .A3(new_n261), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n269), .B1(new_n270), .B2(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n211), .A2(KEYINPUT67), .A3(G20), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT67), .B1(new_n211), .B2(G20), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n229), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n213), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n284), .A2(new_n231), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n287), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n283), .A2(new_n288), .B1(new_n229), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n257), .B1(new_n213), .B2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n212), .B1(new_n228), .B2(new_n229), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n212), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n292), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n279), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n277), .A2(new_n278), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT68), .B1(new_n277), .B2(G169), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n301), .B(KEYINPUT9), .Z(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G200), .B2(new_n276), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n276), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n305), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n282), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n288), .A2(G68), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT77), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n297), .A2(G50), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT76), .Z(new_n320));
  OAI22_X1  g0120(.A1(new_n295), .A2(new_n270), .B1(new_n212), .B2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n292), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n289), .A2(new_n203), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT11), .B(new_n292), .C1(new_n320), .C2(new_n321), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n318), .A2(new_n324), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n267), .A2(new_n268), .ZN(new_n331));
  INV_X1    g0131(.A(G226), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n329), .B1(new_n330), .B2(new_n207), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(new_n274), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n263), .A2(G238), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n265), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT13), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n274), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n328), .B1(G200), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n345), .A2(new_n347), .A3(G190), .A4(new_n341), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n334), .A2(KEYINPUT13), .A3(new_n336), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n350), .B2(new_n346), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n345), .A2(new_n347), .A3(G179), .A4(new_n341), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n342), .A2(new_n354), .A3(G169), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n328), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n295), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G20), .B2(G77), .ZN(new_n360));
  INV_X1    g0160(.A(new_n294), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n291), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n288), .A2(G77), .A3(new_n316), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n289), .A2(new_n270), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g0169(.A(KEYINPUT69), .B(G107), .Z(new_n370));
  OAI22_X1  g0170(.A1(new_n271), .A2(new_n219), .B1(new_n370), .B2(new_n267), .ZN(new_n371));
  INV_X1    g0171(.A(new_n267), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n372), .A2(new_n237), .A3(G1698), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n274), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n263), .A2(G244), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n374), .A2(new_n265), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n369), .B(KEYINPUT72), .C1(G169), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT72), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n375), .A2(new_n265), .ZN(new_n379));
  AOI21_X1  g0179(.A(G169), .B1(new_n379), .B2(new_n374), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n365), .A2(new_n368), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n278), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n379), .B2(new_n374), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT70), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n379), .A2(new_n374), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n386), .A2(new_n387), .B1(new_n388), .B2(new_n308), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n379), .A2(KEYINPUT70), .A3(new_n374), .A4(G190), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(new_n381), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT73), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n393), .A2(KEYINPUT73), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n315), .A2(new_n357), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n204), .A2(new_n205), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G20), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n297), .A2(G159), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n403), .A3(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n267), .B2(G20), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT3), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(G33), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT7), .B(new_n212), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n203), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n397), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n404), .A2(new_n402), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n403), .B1(new_n399), .B2(G20), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(KEYINPUT78), .A3(new_n411), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT78), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n406), .C1(new_n267), .C2(G20), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(G68), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n420), .A3(KEYINPUT16), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n421), .A3(new_n292), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n282), .A2(new_n294), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n288), .B1(new_n289), .B2(new_n294), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n263), .A2(G232), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n408), .A2(G33), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(G226), .A4(G1698), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(G223), .A4(new_n268), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n274), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n425), .A2(new_n434), .A3(new_n308), .A4(new_n265), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n425), .A2(new_n434), .A3(new_n265), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(G200), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n422), .A2(new_n424), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n422), .A2(new_n424), .A3(new_n437), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n439), .B1(new_n444), .B2(KEYINPUT17), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n425), .A2(new_n434), .A3(new_n265), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G169), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(G179), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n422), .A2(new_n424), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT18), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n396), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n208), .A2(KEYINPUT6), .ZN(new_n453));
  OR2_X1    g0253(.A1(KEYINPUT83), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT83), .A2(G97), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G97), .A2(G107), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT6), .B1(new_n209), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G20), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n270), .B2(new_n298), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n370), .B1(new_n407), .B2(new_n411), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n292), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n287), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n211), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n291), .A2(new_n287), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(G97), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n260), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G257), .A3(new_n258), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n258), .A2(G274), .A3(new_n470), .A4(new_n469), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n429), .A2(new_n430), .A3(G250), .A4(G1698), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n429), .A2(new_n430), .A3(G244), .A4(new_n268), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n274), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n477), .A2(G179), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n472), .A2(new_n473), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n274), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n478), .B(KEYINPUT84), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G169), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n468), .B1(G200), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n477), .A2(G190), .A3(new_n487), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n468), .A2(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n504), .B(new_n505), .C1(new_n331), .C2(new_n221), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n274), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n471), .A2(G264), .A3(new_n258), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n473), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n385), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT88), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(KEYINPUT87), .A3(new_n308), .A4(new_n473), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n507), .A2(new_n308), .A3(new_n508), .A4(new_n473), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n509), .A2(KEYINPUT88), .A3(new_n385), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n512), .A2(new_n514), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n267), .A2(new_n212), .A3(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n267), .A2(new_n522), .A3(new_n212), .A4(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT24), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n208), .A2(G20), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  OAI22_X1  g0327(.A1(KEYINPUT23), .A2(new_n526), .B1(new_n295), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n370), .A2(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(KEYINPUT23), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n525), .B1(new_n524), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n292), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n286), .A2(G20), .A3(new_n208), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G107), .B2(new_n466), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n519), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  XOR2_X1   g0340(.A(KEYINPUT83), .B(G97), .Z(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n295), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n267), .A2(new_n212), .A3(G68), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n330), .A2(new_n207), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(new_n545), .B2(KEYINPUT19), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT69), .B(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G87), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n292), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n289), .A2(new_n358), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n466), .A2(G87), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n267), .A2(G238), .A3(new_n268), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n267), .A2(G244), .A3(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n274), .ZN(new_n558));
  AOI21_X1  g0358(.A(G250), .B1(new_n211), .B2(G45), .ZN(new_n559));
  INV_X1    g0359(.A(G274), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n470), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n258), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n558), .A2(G190), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  AOI221_X4 g0366(.A(G179), .B1(new_n258), .B2(new_n561), .C1(new_n557), .C2(new_n274), .ZN(new_n567));
  AOI21_X1  g0367(.A(G169), .B1(new_n558), .B2(new_n562), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n550), .B(new_n551), .C1(new_n358), .C2(new_n465), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n564), .A2(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n503), .A2(new_n539), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n466), .A2(KEYINPUT86), .A3(G116), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n465), .B2(new_n527), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n212), .A2(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n286), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n212), .B(new_n485), .C1(new_n541), .C2(G33), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n291), .A2(new_n578), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT20), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n577), .B(new_n579), .C1(new_n582), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n267), .A2(G257), .A3(new_n268), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  INV_X1    g0387(.A(G264), .ZN(new_n588));
  OAI221_X1 g0388(.A(new_n586), .B1(new_n587), .B2(new_n267), .C1(new_n271), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n274), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n471), .A2(G270), .A3(new_n258), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n591), .A2(new_n473), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n498), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(new_n592), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n278), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n585), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n585), .A2(KEYINPUT21), .A3(new_n593), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n509), .A2(new_n498), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G179), .B2(new_n509), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n538), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n597), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n385), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n597), .A2(new_n308), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n606), .A2(new_n607), .A3(new_n585), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n601), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n452), .A2(new_n573), .A3(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n356), .A2(new_n328), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n349), .B2(new_n384), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n445), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n450), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n312), .A2(new_n314), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n305), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n452), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT89), .ZN(new_n618));
  INV_X1    g0418(.A(new_n488), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n498), .B1(new_n477), .B2(new_n487), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n468), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n468), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n622), .B(new_n502), .C1(new_n497), .C2(new_n385), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n571), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n509), .A2(KEYINPUT88), .A3(new_n385), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT88), .B1(new_n509), .B2(new_n385), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n515), .B(KEYINPUT87), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n537), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n618), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n503), .A2(new_n539), .A3(KEYINPUT89), .A4(new_n571), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n537), .B(new_n602), .C1(G179), .C2(new_n509), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n596), .A3(new_n599), .A4(new_n600), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n553), .ZN(new_n635));
  INV_X1    g0435(.A(new_n563), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n566), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n569), .A2(new_n570), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n499), .A2(new_n637), .A3(new_n638), .A4(new_n468), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .B1(new_n570), .B2(new_n569), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n622), .B1(new_n499), .B2(KEYINPUT90), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n488), .B(new_n643), .C1(new_n497), .C2(new_n498), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n571), .A4(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n616), .B1(new_n617), .B2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n286), .A2(new_n212), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT91), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  AND4_X1   g0453(.A1(G213), .A2(new_n652), .A3(G343), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n585), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n601), .B(new_n655), .Z(new_n656));
  INV_X1    g0456(.A(new_n608), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(KEYINPUT92), .B(G330), .Z(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n654), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n538), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n632), .B1(new_n629), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n604), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n664), .A2(new_n601), .A3(new_n632), .A4(new_n662), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n665), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n215), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n230), .ZN(new_n674));
  OAI21_X1  g0474(.A(G1), .B1(new_n672), .B2(G41), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n548), .A2(new_n527), .A3(new_n541), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(new_n639), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n679), .A2(new_n642), .B1(new_n570), .B2(new_n569), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n641), .A2(new_n571), .A3(new_n644), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n682));
  INV_X1    g0482(.A(new_n633), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n680), .B(new_n682), .C1(new_n572), .C2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(KEYINPUT29), .A3(new_n662), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n654), .B1(new_n634), .B2(new_n646), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(KEYINPUT29), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n573), .A2(new_n609), .A3(new_n662), .ZN(new_n688));
  AND4_X1   g0488(.A1(new_n508), .A2(new_n507), .A3(new_n562), .A4(new_n558), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n598), .A2(new_n497), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n605), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n509), .A3(new_n565), .A4(new_n500), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n598), .A2(new_n497), .A3(KEYINPUT30), .A4(new_n689), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n654), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n688), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n659), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n687), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n678), .B1(new_n704), .B2(G1), .ZN(G364));
  NOR2_X1   g0505(.A1(new_n285), .A2(G20), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n211), .B1(new_n706), .B2(G45), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OR3_X1    g0508(.A1(new_n673), .A2(KEYINPUT93), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT93), .B1(new_n673), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n658), .A2(new_n659), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n661), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G13), .A2(G33), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n658), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n212), .A2(G179), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n308), .A3(G200), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n721));
  OAI221_X1 g0521(.A(new_n267), .B1(new_n720), .B2(new_n208), .C1(new_n220), .C2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n212), .A2(new_n278), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT97), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT97), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n308), .A2(G200), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G190), .A2(G200), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n202), .A2(new_n727), .B1(new_n729), .B2(new_n270), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n723), .A2(G190), .A3(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT98), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n731), .A2(KEYINPUT98), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n722), .B(new_n730), .C1(G50), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n719), .A2(new_n728), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT99), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT99), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G159), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT32), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n212), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n207), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n723), .A2(new_n308), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(G68), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT100), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n737), .A2(new_n744), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(KEYINPUT33), .A2(G317), .ZN(new_n753));
  AND2_X1   g0553(.A1(KEYINPUT33), .A2(G317), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n755), .B1(new_n756), .B2(new_n746), .C1(new_n587), .C2(new_n721), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(G326), .B2(new_n736), .ZN(new_n758));
  INV_X1    g0558(.A(new_n727), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G322), .ZN(new_n760));
  INV_X1    g0560(.A(new_n720), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n267), .B1(new_n761), .B2(G283), .ZN(new_n762));
  INV_X1    g0562(.A(new_n741), .ZN(new_n763));
  INV_X1    g0563(.A(new_n729), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(G329), .B1(new_n764), .B2(G311), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n758), .A2(new_n760), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n752), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n231), .B1(G20), .B2(new_n498), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n711), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n672), .A2(new_n372), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G355), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G116), .B2(new_n215), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n251), .A2(G45), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT95), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n672), .A2(new_n267), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n230), .B2(new_n260), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n772), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(KEYINPUT96), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT96), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n717), .A2(new_n768), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n718), .B(new_n769), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n714), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT101), .Z(G396));
  INV_X1    g0585(.A(new_n711), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT103), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n654), .A2(new_n369), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n384), .A2(new_n787), .A3(new_n392), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n788), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n790), .A2(new_n382), .A3(new_n383), .A4(new_n377), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n384), .A2(new_n392), .A3(new_n788), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT103), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n686), .B(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n786), .B1(new_n796), .B2(new_n703), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n703), .B2(new_n796), .ZN(new_n798));
  INV_X1    g0598(.A(new_n768), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n716), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n786), .B1(G77), .B2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n763), .A2(G311), .B1(G87), .B2(new_n761), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT102), .Z(new_n803));
  OAI22_X1  g0603(.A1(new_n527), .A2(new_n729), .B1(new_n727), .B2(new_n756), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n748), .A2(new_n805), .B1(new_n721), .B2(new_n208), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n804), .A2(new_n267), .A3(new_n747), .A4(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n803), .B(new_n807), .C1(new_n587), .C2(new_n735), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n759), .A2(G143), .B1(G150), .B2(new_n749), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n742), .B2(new_n729), .C1(new_n810), .C2(new_n735), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  INV_X1    g0612(.A(new_n721), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G50), .B1(new_n761), .B2(G68), .ZN(new_n814));
  INV_X1    g0614(.A(new_n746), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n372), .B1(new_n815), .B2(G58), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n814), .B(new_n816), .C1(new_n741), .C2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n808), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n801), .B1(new_n819), .B2(new_n768), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n795), .B2(new_n716), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n798), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  OR2_X1    g0623(.A1(new_n456), .A2(new_n458), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT35), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(KEYINPUT35), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n825), .A2(G116), .A3(new_n232), .A4(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  NAND3_X1  g0628(.A1(new_n230), .A2(G77), .A3(new_n398), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n229), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n211), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT104), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n647), .A2(new_n662), .A3(new_n795), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n384), .A2(new_n654), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n343), .A2(new_n348), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n328), .A2(new_n654), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n611), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n328), .B(new_n654), .C1(new_n349), .C2(new_n356), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n833), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n421), .A2(new_n292), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n416), .A2(new_n420), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n397), .ZN(new_n848));
  INV_X1    g0648(.A(new_n424), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n445), .B2(new_n450), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n444), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n422), .A2(new_n424), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n851), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n858), .A2(KEYINPUT37), .A3(new_n449), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n448), .A2(new_n447), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n848), .A2(new_n849), .B1(new_n860), .B2(new_n851), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n441), .A3(new_n443), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n855), .A2(new_n859), .B1(new_n862), .B2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n853), .B2(new_n863), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n837), .A2(KEYINPUT104), .A3(new_n843), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n845), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n450), .A2(new_n851), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  XOR2_X1   g0673(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n438), .B2(new_n449), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n856), .A2(new_n860), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(KEYINPUT106), .A3(new_n442), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n878), .A3(new_n857), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n855), .A2(new_n859), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n451), .A2(new_n858), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n874), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n853), .A2(new_n866), .A3(new_n863), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n611), .A2(new_n654), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n865), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n872), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n452), .B(new_n685), .C1(KEYINPUT29), .C2(new_n686), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n616), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n893), .B(new_n895), .Z(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT108), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n887), .B2(new_n888), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n880), .A2(new_n881), .B1(new_n855), .B2(new_n859), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n900), .A2(new_n884), .B1(new_n451), .B2(new_n858), .ZN(new_n901));
  OAI211_X1 g0701(.A(KEYINPUT108), .B(new_n865), .C1(new_n901), .C2(new_n874), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n841), .A2(new_n842), .B1(new_n792), .B2(new_n794), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n701), .A2(new_n903), .A3(KEYINPUT40), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n899), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n701), .A2(new_n903), .ZN(new_n906));
  INV_X1    g0706(.A(new_n867), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n907), .B2(new_n888), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n452), .A2(new_n701), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n914), .A2(new_n915), .A3(new_n659), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n897), .A2(new_n916), .B1(new_n211), .B2(new_n706), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n897), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n832), .B1(new_n917), .B2(new_n918), .ZN(G367));
  OAI21_X1  g0719(.A(new_n571), .B1(new_n635), .B2(new_n662), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n654), .A2(new_n569), .A3(new_n570), .A4(new_n553), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n503), .B1(new_n622), .B2(new_n662), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n641), .A2(new_n644), .A3(new_n654), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(new_n669), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n926), .A2(new_n604), .B1(new_n468), .B2(new_n499), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n654), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n668), .A2(new_n927), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n673), .B(KEYINPUT41), .Z(new_n938));
  NOR2_X1   g0738(.A1(new_n670), .A2(new_n926), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT44), .Z(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n670), .B2(new_n926), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n670), .A2(new_n941), .A3(new_n926), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT45), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n668), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n601), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n666), .B1(new_n950), .B2(new_n654), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n669), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n660), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n704), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n668), .B1(new_n946), .B2(new_n947), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n938), .B1(new_n956), .B2(new_n704), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n937), .B1(new_n957), .B2(new_n708), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n781), .B1(new_n215), .B2(new_n358), .C1(new_n776), .C2(new_n243), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n960), .A2(new_n961), .A3(new_n711), .ZN(new_n962));
  INV_X1    g0762(.A(new_n717), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G68), .A2(new_n815), .B1(new_n749), .B2(G159), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n720), .A2(new_n270), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(new_n372), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n964), .B1(new_n202), .B2(new_n721), .C1(KEYINPUT112), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n968));
  INV_X1    g0768(.A(G143), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n735), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G50), .A2(new_n764), .B1(new_n759), .B2(G150), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n810), .C2(new_n741), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n813), .A2(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n729), .A2(new_n805), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n746), .A2(new_n370), .B1(new_n541), .B2(new_n720), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n267), .B(new_n978), .C1(G294), .C2(new_n749), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n736), .A2(G311), .ZN(new_n980));
  XNOR2_X1  g0780(.A(KEYINPUT111), .B(G317), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n763), .A2(new_n982), .B1(new_n759), .B2(G303), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n962), .B1(new_n963), .B2(new_n922), .C1(new_n987), .C2(new_n799), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n958), .A2(new_n988), .ZN(G387));
  OR2_X1    g0789(.A1(new_n240), .A2(new_n260), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n990), .A2(new_n775), .B1(new_n676), .B2(new_n770), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n294), .A2(G50), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT50), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n260), .B1(new_n203), .B2(new_n270), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n676), .B(new_n994), .C1(new_n993), .C2(new_n992), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n991), .A2(new_n995), .B1(G107), .B2(new_n215), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n711), .B1(new_n996), .B2(new_n781), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n746), .A2(new_n358), .B1(new_n748), .B2(new_n294), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n759), .B2(G50), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n736), .A2(KEYINPUT115), .A3(G159), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT115), .B1(new_n736), .B2(G159), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n999), .B1(new_n203), .B2(new_n729), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n813), .A2(G77), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n372), .B1(new_n761), .B2(G97), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n741), .C2(new_n296), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT114), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n372), .B1(new_n720), .B2(new_n527), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n764), .A2(G303), .B1(G311), .B2(new_n749), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT116), .B(G322), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n727), .B2(new_n981), .C1(new_n735), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n815), .A2(G283), .B1(new_n813), .B2(G294), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1008), .B(new_n1018), .C1(G326), .C2(new_n763), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1007), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n997), .B1(new_n1021), .B2(new_n799), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n666), .B2(new_n717), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n953), .B2(new_n708), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n673), .B(KEYINPUT117), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n954), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n953), .A2(new_n704), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(G393));
  OAI21_X1  g0828(.A(new_n954), .B1(new_n949), .B2(new_n955), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n956), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n949), .A2(new_n707), .A3(new_n955), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n927), .A2(new_n717), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n248), .A2(new_n775), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n781), .B1(new_n215), .B2(new_n541), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n786), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n736), .A2(G317), .B1(new_n759), .B2(G311), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G116), .A2(new_n815), .B1(new_n749), .B2(G303), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n805), .B2(new_n721), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n267), .B1(new_n761), .B2(G107), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n729), .B2(new_n756), .C1(new_n741), .C2(new_n1010), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n735), .A2(new_n296), .B1(new_n742), .B2(new_n727), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT51), .Z(new_n1044));
  AOI22_X1  g0844(.A1(G50), .A2(new_n749), .B1(new_n813), .B2(G68), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n270), .B2(new_n746), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n372), .B1(new_n761), .B2(G87), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n729), .B2(new_n294), .C1(new_n741), .C2(new_n969), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1035), .B1(new_n1050), .B2(new_n768), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1031), .B1(new_n1032), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1030), .A2(new_n1052), .ZN(G390));
  INV_X1    g0853(.A(G330), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n699), .A2(new_n700), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n688), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n903), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n684), .A2(new_n795), .A3(new_n662), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n836), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n890), .B1(new_n1060), .B2(new_n843), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n899), .A2(new_n902), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n890), .B1(new_n837), .B2(new_n843), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n889), .B2(new_n891), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1058), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT118), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n701), .A2(new_n702), .A3(new_n795), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(new_n844), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT118), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n1058), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1056), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n894), .B(new_n616), .C1(new_n617), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1068), .A2(new_n844), .ZN(new_n1075));
  OAI211_X1 g0875(.A(KEYINPUT119), .B(new_n837), .C1(new_n1075), .C2(new_n1058), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT119), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1068), .A2(new_n844), .B1(new_n1056), .B2(new_n903), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n838), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n795), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n844), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1082), .A2(new_n1069), .A3(new_n836), .A4(new_n1059), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1074), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1066), .A2(new_n1070), .A3(new_n1072), .A4(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1085), .A2(new_n1025), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1066), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1084), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1066), .A2(new_n1070), .A3(new_n708), .A4(new_n1072), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n815), .A2(G77), .B1(new_n761), .B2(G68), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n370), .B2(new_n748), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n729), .A2(new_n541), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n267), .B1(new_n813), .B2(G87), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n527), .B2(new_n727), .C1(new_n756), .C2(new_n741), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1093), .B(new_n1097), .C1(G283), .C2(new_n736), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n721), .A2(new_n296), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G125), .B2(new_n763), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n817), .A2(new_n727), .B1(new_n729), .B2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n748), .A2(new_n810), .B1(new_n720), .B2(new_n229), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n372), .B(new_n1105), .C1(G159), .C2(new_n815), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(G128), .C2(new_n736), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1098), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n786), .B1(new_n361), .B2(new_n800), .C1(new_n1109), .C2(new_n799), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n889), .A2(new_n891), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n716), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1091), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1090), .A2(new_n1115), .ZN(G378));
  AOI21_X1  g0916(.A(new_n1054), .B1(new_n908), .B2(new_n909), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n905), .A2(new_n1117), .A3(KEYINPUT122), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT122), .B1(new_n905), .B2(new_n1117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n851), .A2(new_n301), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n315), .B(new_n1120), .Z(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1124), .A2(KEYINPUT122), .A3(new_n905), .A4(new_n1117), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1125), .A2(new_n1127), .B1(new_n892), .B2(new_n872), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n905), .A2(new_n1117), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT122), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n905), .A2(new_n1117), .A3(KEYINPUT122), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1123), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n893), .A3(new_n1126), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n708), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n786), .B1(G50), .B2(new_n800), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n267), .A2(G41), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G50), .B(new_n1137), .C1(new_n330), .C2(new_n259), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1137), .B1(new_n203), .B2(new_n746), .C1(new_n741), .C2(new_n805), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n735), .A2(new_n527), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n208), .A2(new_n727), .B1(new_n729), .B2(new_n358), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1003), .B1(new_n202), .B2(new_n720), .C1(new_n207), .C2(new_n748), .ZN(new_n1142));
  OR4_X1    g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT58), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1138), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n736), .A2(G125), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G128), .A2(new_n759), .B1(new_n764), .B2(G137), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1103), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n813), .A2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G150), .A2(new_n815), .B1(new_n749), .B2(G132), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n763), .A2(G124), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G33), .B(G41), .C1(new_n761), .C2(G159), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1145), .B1(new_n1144), .B2(new_n1143), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1136), .B1(new_n1157), .B2(new_n768), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1123), .B2(new_n716), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT121), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1135), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1074), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1085), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(KEYINPUT57), .A3(new_n1134), .A4(new_n1128), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1025), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1133), .A2(new_n893), .A3(new_n1126), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n893), .B1(new_n1133), .B2(new_n1126), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1163), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1161), .B1(new_n1165), .B2(new_n1169), .ZN(G375));
  NAND2_X1  g0970(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n844), .A2(new_n715), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n786), .B1(G68), .B2(new_n800), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n267), .B(new_n965), .C1(new_n763), .C2(G303), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n805), .B2(new_n727), .C1(new_n370), .C2(new_n729), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n358), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1176), .A2(new_n815), .B1(new_n749), .B2(G116), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n207), .B2(new_n721), .C1(new_n735), .C2(new_n756), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n267), .B1(new_n720), .B2(new_n202), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n763), .B2(G128), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n810), .B2(new_n727), .C1(new_n296), .C2(new_n729), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G50), .A2(new_n815), .B1(new_n749), .B2(new_n1148), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n742), .B2(new_n721), .C1(new_n735), .C2(new_n817), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1175), .A2(new_n1178), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1173), .B1(new_n1184), .B2(new_n768), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1171), .A2(new_n708), .B1(new_n1172), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n938), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1088), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1171), .A2(new_n1162), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(G381));
  OR2_X1    g0990(.A1(G375), .A2(G378), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n784), .B(KEYINPUT101), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1024), .C1(new_n1027), .C2(new_n1026), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1194), .A2(new_n822), .A3(new_n1030), .A4(new_n1052), .ZN(new_n1195));
  OR4_X1    g0995(.A1(G387), .A2(new_n1191), .A3(G381), .A4(new_n1195), .ZN(G407));
  OAI211_X1 g0996(.A(G407), .B(G213), .C1(G343), .C2(new_n1191), .ZN(G409));
  AND2_X1   g0997(.A1(G396), .A2(G393), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(G390), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1052), .B(new_n1030), .C1(new_n1194), .C2(new_n1198), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(G387), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT61), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1200), .A2(new_n1201), .A3(new_n958), .A4(new_n988), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G378), .B(new_n1161), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1114), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1168), .A2(new_n1187), .A3(new_n1163), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1135), .A2(new_n1160), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(G343), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(G213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1171), .B2(new_n1162), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1215), .A2(new_n1025), .A3(new_n1088), .A4(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(G384), .A3(new_n1186), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G384), .B1(new_n1218), .B2(new_n1186), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1212), .A2(new_n1214), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1206), .B1(new_n1224), .B2(KEYINPUT63), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1214), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(G2897), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT125), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n1222), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1229), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1227), .A2(KEYINPUT124), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(KEYINPUT124), .B2(new_n1227), .ZN(new_n1234));
  AOI211_X1 g1034(.A(KEYINPUT123), .B(KEYINPUT63), .C1(new_n1227), .C2(new_n1222), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT123), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1223), .B2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1225), .B(new_n1234), .C1(new_n1235), .C2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1227), .A2(KEYINPUT62), .A3(new_n1222), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT62), .B1(new_n1227), .B2(new_n1222), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1242), .B(KEYINPUT126), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1223), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1227), .A2(KEYINPUT62), .A3(new_n1222), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT126), .B1(new_n1251), .B2(new_n1242), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1239), .B1(new_n1247), .B2(new_n1252), .ZN(G405));
  INV_X1    g1053(.A(KEYINPUT127), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1222), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1246), .B(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1222), .A2(new_n1254), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1207), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1208), .B2(G375), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1256), .B(new_n1259), .ZN(G402));
endmodule


