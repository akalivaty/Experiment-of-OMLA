//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT24), .B(G110), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n197), .B2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  INV_X1    g020(.A(G110), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n198), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n209), .A2(KEYINPUT74), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(KEYINPUT74), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n193), .B(new_n196), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n196), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n206), .A3(new_n198), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G110), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT73), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n201), .A2(new_n202), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n215), .B(new_n217), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n224), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT75), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n212), .A2(new_n222), .A3(KEYINPUT75), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n227), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G234), .ZN(new_n236));
  OAI21_X1  g050(.A(G217), .B1(new_n236), .B2(G902), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n235), .B2(G902), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n212), .A2(new_n222), .A3(KEYINPUT75), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT75), .B1(new_n212), .B2(new_n222), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n234), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n228), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n237), .B(KEYINPUT72), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n242), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT66), .A2(G134), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT66), .A2(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n263), .B1(G134), .B2(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(G128), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n192), .A2(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(G146), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(new_n265), .B2(G146), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n192), .A3(G143), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n270), .A4(new_n276), .ZN(new_n277));
  AOI22_X1  g091(.A1(G131), .A2(new_n264), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n260), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n263), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n261), .A2(new_n262), .ZN(new_n283));
  AOI21_X1  g097(.A(G131), .B1(new_n283), .B2(G137), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT67), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g101(.A1(KEYINPUT2), .A2(G113), .ZN(new_n288));
  AND3_X1   g102(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n197), .A2(G116), .ZN(new_n292));
  INV_X1    g106(.A(G116), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G119), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G116), .B(G119), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n288), .C1(new_n290), .C2(new_n289), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT69), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(new_n300), .A3(new_n295), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n283), .A2(G137), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n282), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n306));
  OR2_X1    g120(.A1(KEYINPUT66), .A2(G134), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT66), .A2(G134), .ZN(new_n308));
  AOI21_X1  g122(.A(G137), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n279), .B1(new_n309), .B2(KEYINPUT11), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n303), .B1(new_n311), .B2(new_n260), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n284), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n305), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT0), .A2(G128), .ZN(new_n316));
  OR2_X1    g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n271), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n273), .A2(new_n275), .A3(new_n270), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n287), .B(new_n302), .C1(new_n315), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n302), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n313), .A2(new_n314), .ZN(new_n325));
  INV_X1    g139(.A(new_n304), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n310), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n287), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n278), .C1(new_n285), .C2(new_n286), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n325), .B2(new_n278), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n327), .B1(new_n285), .B2(new_n286), .ZN(new_n337));
  INV_X1    g151(.A(new_n320), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n336), .A2(KEYINPUT28), .A3(new_n302), .A4(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n259), .B1(new_n331), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT30), .A4(new_n333), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n328), .B2(new_n329), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n344), .A2(new_n324), .A3(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n339), .A2(new_n343), .A3(new_n302), .A4(new_n333), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n259), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n342), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(new_n346), .A3(new_n324), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT31), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n341), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(G472), .A2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n348), .A2(new_n322), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n323), .A2(new_n330), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n259), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n259), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n352), .A2(new_n361), .A3(new_n348), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n323), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n339), .A2(new_n343), .A3(new_n333), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n324), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n348), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n361), .A2(new_n364), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(KEYINPUT32), .A2(new_n357), .B1(new_n373), .B2(G472), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n354), .B2(new_n356), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n361), .B1(new_n358), .B2(new_n359), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n347), .A2(new_n342), .A3(new_n349), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT31), .B1(new_n351), .B2(new_n352), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT71), .A3(new_n355), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT32), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n254), .B1(new_n374), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G116), .B(G122), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n265), .A2(G128), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT13), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n199), .A2(G143), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  OAI21_X1  g207(.A(G134), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n391), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n387), .B(new_n394), .C1(new_n311), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n293), .A3(G122), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n293), .B2(G122), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n293), .B2(G122), .ZN(new_n400));
  OAI21_X1  g214(.A(G107), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT97), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n311), .B(new_n395), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n386), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n396), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT9), .B(G234), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(G217), .A3(new_n225), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n406), .A2(new_n409), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G902), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G237), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(new_n225), .A3(G143), .A4(G214), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n255), .A2(new_n421), .A3(G143), .A4(G214), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G214), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(G237), .A3(G953), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n425), .A2(new_n426), .A3(G143), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n255), .A2(G214), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT88), .B1(new_n428), .B2(new_n265), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n423), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(KEYINPUT18), .A2(G131), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n191), .A2(new_n192), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT91), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n193), .A2(KEYINPUT90), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n426), .B1(new_n425), .B2(G143), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n428), .A2(KEYINPUT88), .A3(new_n265), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n439), .A2(new_n440), .B1(new_n420), .B2(new_n422), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT92), .B1(new_n441), .B2(new_n303), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT92), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n430), .A2(new_n443), .A3(G131), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n214), .A2(KEYINPUT95), .A3(new_n196), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT95), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n215), .A2(new_n447), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n445), .A2(KEYINPUT17), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n441), .A2(new_n303), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n442), .A2(new_n444), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT96), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n452), .A2(new_n453), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n438), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(G104), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n460), .B(new_n438), .C1(new_n455), .C2(new_n456), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G475), .B1(new_n464), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n445), .B1(new_n303), .B2(new_n441), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n191), .A2(KEYINPUT93), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT19), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT94), .B1(new_n469), .B2(G146), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n468), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT94), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n192), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n196), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n438), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n461), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n479), .ZN(new_n481));
  AOI211_X1 g295(.A(KEYINPUT20), .B(new_n481), .C1(new_n477), .C2(new_n463), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n417), .B(new_n465), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n320), .A2(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n272), .A2(new_n277), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(G125), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G224), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(G953), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT84), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n486), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G101), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n386), .A2(G104), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n459), .A2(G107), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT3), .B1(new_n459), .B2(G107), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n386), .A3(G104), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n495), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT80), .B(G101), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g315(.A(G113), .B1(new_n292), .B2(KEYINPUT5), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n500), .B(new_n298), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n499), .A2(new_n495), .A3(new_n493), .A4(new_n497), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n497), .A3(new_n493), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n504), .A2(KEYINPUT4), .B1(G101), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n505), .A2(KEYINPUT4), .A3(G101), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n503), .B1(new_n508), .B2(new_n302), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT83), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n503), .B(KEYINPUT83), .C1(new_n508), .C2(new_n302), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G122), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n511), .A2(KEYINPUT6), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n509), .A2(new_n514), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT6), .B1(new_n519), .B2(new_n512), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n490), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT7), .B1(new_n487), .B2(G953), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n486), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n492), .A2(new_n493), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G101), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n504), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n501), .A2(KEYINPUT85), .ZN(new_n527));
  AND4_X1   g341(.A1(KEYINPUT85), .A2(new_n292), .A3(new_n294), .A4(KEYINPUT5), .ZN(new_n528));
  OR3_X1    g342(.A1(new_n527), .A2(new_n528), .A3(new_n502), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n526), .B1(new_n529), .B2(new_n298), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n513), .B(KEYINPUT8), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n298), .B1(new_n501), .B2(new_n502), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n500), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n523), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n516), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n486), .A2(new_n522), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT86), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n521), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G210), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n521), .A2(new_n538), .A3(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n540), .B1(new_n521), .B2(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(G234), .A2(G237), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(G952), .A3(new_n225), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT21), .B(G898), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(G902), .A3(G953), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n483), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G469), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  INV_X1    g373(.A(G227), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(G953), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n559), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n319), .A2(new_n268), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n277), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n500), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT10), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n338), .B1(new_n506), .B2(new_n507), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n500), .A2(new_n485), .A3(KEYINPUT10), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n315), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n526), .A2(new_n272), .A3(new_n277), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n337), .A2(KEYINPUT12), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT12), .B1(new_n337), .B2(new_n572), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT81), .B(new_n570), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n565), .A2(new_n571), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(new_n315), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n337), .A2(KEYINPUT12), .A3(new_n572), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT81), .B1(new_n581), .B2(new_n570), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n562), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n562), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n570), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n337), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n558), .B1(new_n590), .B2(new_n238), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n581), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n570), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n562), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT82), .B(G469), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n408), .A2(new_n238), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G221), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT79), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n384), .A2(new_n557), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT98), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(new_n499), .Z(G3));
  INV_X1    g420(.A(new_n602), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n253), .B(new_n607), .C1(new_n591), .C2(new_n598), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n354), .B2(G902), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n376), .A2(new_n609), .A3(new_n381), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n521), .A2(new_n538), .A3(new_n540), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n555), .B1(new_n612), .B2(new_n545), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(new_n555), .C1(new_n612), .C2(new_n545), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n614), .A2(new_n554), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n462), .B2(new_n463), .ZN(new_n618));
  INV_X1    g432(.A(G475), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n480), .A2(new_n482), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n413), .A2(new_n414), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n414), .A2(new_n238), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n412), .B(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(G478), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n611), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  OAI211_X1 g445(.A(new_n465), .B(new_n416), .C1(new_n480), .C2(new_n482), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n611), .A2(new_n617), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n386), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(new_n589), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT81), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n575), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n638), .B1(new_n642), .B2(new_n562), .ZN(new_n643));
  OAI21_X1  g457(.A(G469), .B1(new_n643), .B2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n597), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT25), .B1(new_n248), .B2(new_n238), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n243), .B(G902), .C1(new_n247), .C2(new_n228), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n252), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n234), .A2(KEYINPUT36), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n233), .B(new_n649), .Z(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n648), .B1(new_n241), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n645), .A2(new_n607), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n610), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n557), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AOI21_X1  g471(.A(new_n653), .B1(new_n383), .B2(new_n374), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n614), .A2(new_n616), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT101), .B(G900), .Z(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(new_n553), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n550), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n632), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(new_n548), .B(KEYINPUT38), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n380), .A2(KEYINPUT32), .A3(new_n355), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n238), .B1(new_n369), .B2(new_n259), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n361), .B1(new_n352), .B2(new_n348), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(KEYINPUT102), .B(G472), .C1(new_n670), .C2(new_n671), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n669), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n676), .A2(new_n383), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n668), .A2(new_n677), .A3(new_n652), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n620), .A2(new_n416), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n555), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n663), .B(KEYINPUT39), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n603), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n680), .B1(new_n682), .B2(KEYINPUT40), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n678), .B(new_n683), .C1(KEYINPUT40), .C2(new_n682), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND3_X1  g499(.A1(new_n620), .A2(new_n626), .A3(new_n663), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n660), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NOR2_X1   g503(.A1(new_n595), .A2(new_n558), .ZN(new_n690));
  INV_X1    g504(.A(new_n601), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n598), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n384), .A2(new_n617), .A3(new_n628), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND4_X1  g509(.A1(new_n384), .A2(new_n617), .A3(new_n633), .A4(new_n692), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT103), .B(G116), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G18));
  AOI21_X1  g512(.A(new_n483), .B1(new_n374), .B2(new_n383), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n692), .A2(new_n652), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n617), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n302), .B1(new_n336), .B2(new_n339), .ZN(new_n704));
  INV_X1    g518(.A(new_n348), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT28), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n323), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n361), .B1(new_n350), .B2(new_n353), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n703), .B1(new_n708), .B2(new_n356), .ZN(new_n709));
  OAI22_X1  g523(.A1(new_n378), .A2(new_n379), .B1(new_n370), .B2(new_n259), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n355), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n253), .A2(new_n709), .A3(new_n609), .A4(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n617), .A2(new_n712), .A3(new_n679), .A4(new_n692), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NAND2_X1  g528(.A1(new_n710), .A2(new_n355), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n380), .A2(new_n238), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n703), .A2(new_n715), .B1(new_n716), .B2(G472), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n687), .A2(new_n652), .A3(new_n717), .A4(new_n711), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n614), .A2(new_n616), .A3(new_n692), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n709), .A2(new_n609), .A3(new_n652), .A4(new_n711), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n686), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  INV_X1    g537(.A(new_n719), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND2_X1  g541(.A1(new_n373), .A2(G472), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n382), .B1(new_n354), .B2(new_n356), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n669), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n687), .A2(new_n253), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n555), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n544), .B2(new_n547), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n691), .B1(new_n644), .B2(new_n597), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT42), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n548), .A2(new_n734), .A3(new_n555), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n384), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n303), .ZN(G33));
  NAND2_X1  g555(.A1(new_n374), .A2(new_n383), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n742), .A3(new_n253), .A4(new_n665), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n384), .A2(new_n737), .A3(KEYINPUT106), .A4(new_n665), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NAND2_X1  g562(.A1(new_n625), .A2(G478), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n621), .A3(new_n623), .ZN(new_n750));
  OR3_X1    g564(.A1(new_n620), .A2(new_n750), .A3(KEYINPUT43), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT43), .B1(new_n620), .B2(new_n750), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n610), .A3(new_n652), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT107), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n643), .A2(KEYINPUT45), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n643), .A2(KEYINPUT45), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(G469), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(G469), .A2(G902), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT46), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n598), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n760), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n691), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n681), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n733), .B1(new_n753), .B2(new_n754), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n756), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  OR2_X1    g582(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n733), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n742), .A2(new_n772), .A3(new_n253), .A4(new_n686), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT108), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(new_n712), .ZN(new_n777));
  INV_X1    g591(.A(new_n550), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n751), .A2(new_n778), .A3(new_n752), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n668), .A2(new_n732), .A3(new_n692), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n781), .A2(new_n782), .ZN(new_n788));
  INV_X1    g602(.A(new_n721), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n733), .A2(new_n692), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT115), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n788), .A2(new_n793), .A3(new_n789), .A4(new_n790), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n778), .A2(new_n677), .A3(new_n253), .A4(new_n790), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n620), .A2(new_n626), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n792), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n783), .A2(new_n733), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n764), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n598), .A2(new_n690), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n602), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n798), .A2(KEYINPUT116), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n787), .A2(new_n797), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n769), .A2(new_n809), .A3(new_n770), .A4(new_n803), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n799), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n801), .B2(new_n803), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT51), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n787), .A4(new_n797), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT118), .B1(new_n798), .B2(new_n813), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n795), .A2(new_n628), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(G952), .A3(new_n225), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n783), .B2(new_n724), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n730), .A2(new_n253), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n788), .A2(new_n822), .A3(new_n790), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT48), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT119), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(KEYINPUT119), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n823), .A2(new_n826), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n820), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT120), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n820), .A2(new_n829), .A3(new_n832), .A4(new_n828), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n816), .A2(new_n817), .A3(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n808), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n772), .A2(new_n653), .A3(new_n664), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n699), .B1(new_n722), .B2(new_n737), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n747), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n747), .A2(KEYINPUT111), .A3(new_n838), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n548), .A2(new_n556), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n632), .B2(new_n627), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT110), .B1(new_n620), .B2(new_n626), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n611), .B(new_n843), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n693), .A2(new_n696), .A3(new_n847), .A4(new_n701), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n713), .A2(new_n604), .A3(new_n655), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n848), .A2(new_n740), .A3(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n841), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n658), .B(new_n659), .C1(new_n665), .C2(new_n687), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n652), .B1(new_n676), .B2(new_n383), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n734), .A2(new_n663), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n659), .A3(new_n679), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n723), .B1(new_n722), .B2(new_n724), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n719), .A2(new_n721), .A3(KEYINPUT105), .A4(new_n686), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n852), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n726), .A2(KEYINPUT52), .A3(new_n852), .A4(new_n855), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT112), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n851), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n841), .A2(new_n842), .A3(new_n850), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n860), .A2(new_n861), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT54), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT113), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n873), .B(new_n865), .C1(new_n867), .C2(new_n868), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n851), .B(KEYINPUT53), .C1(new_n862), .C2(new_n863), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(KEYINPUT54), .B2(new_n876), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n836), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  INV_X1    g692(.A(new_n802), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(KEYINPUT49), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT109), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(KEYINPUT49), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n555), .A3(new_n253), .A4(new_n607), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n881), .A2(new_n620), .A3(new_n750), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n677), .A3(new_n668), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n878), .A2(new_n885), .ZN(G75));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n876), .A2(G902), .ZN(new_n888));
  INV_X1    g702(.A(G210), .ZN(new_n889));
  OAI211_X1 g703(.A(KEYINPUT122), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n518), .A2(new_n520), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT121), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n490), .B(KEYINPUT55), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n225), .A2(G952), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n890), .B2(new_n894), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n592), .A2(new_n594), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n876), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n760), .B(KEYINPUT57), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n888), .A2(new_n759), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n896), .B1(new_n904), .B2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n907));
  INV_X1    g721(.A(new_n478), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n896), .ZN(G60));
  XOR2_X1   g725(.A(new_n625), .B(KEYINPUT123), .Z(new_n912));
  XOR2_X1   g726(.A(new_n622), .B(KEYINPUT59), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n897), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n877), .B2(new_n913), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  NAND3_X1  g733(.A1(new_n876), .A2(new_n650), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n876), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n235), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n876), .A2(KEYINPUT125), .A3(new_n650), .A4(new_n919), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n924), .A3(new_n897), .A4(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n897), .A4(new_n920), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  NOR2_X1   g744(.A1(new_n848), .A2(new_n849), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n225), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT126), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n551), .B2(new_n487), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(G898), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n892), .B1(new_n937), .B2(G953), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n936), .B(new_n938), .Z(G69));
  NAND3_X1  g753(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n344), .A2(new_n346), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n469), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n684), .A2(new_n726), .A3(new_n852), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  NOR2_X1   g759(.A1(new_n682), .A2(new_n772), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n384), .C1(new_n845), .C2(new_n846), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n945), .A2(new_n775), .A3(new_n767), .A4(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n940), .B(new_n943), .C1(new_n948), .C2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n726), .A2(new_n852), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n822), .A2(new_n659), .A3(new_n679), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n765), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n747), .ZN(new_n953));
  NOR4_X1   g767(.A1(new_n950), .A2(new_n952), .A3(new_n953), .A4(new_n740), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n775), .A2(new_n767), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(G953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n560), .A2(G900), .A3(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n942), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n949), .B1(new_n959), .B2(new_n961), .ZN(G72));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n931), .A3(new_n958), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  AOI21_X1  g779(.A(new_n362), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n948), .B2(new_n932), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n671), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n897), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n866), .A2(new_n869), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n362), .A2(new_n965), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n970), .A2(new_n671), .A3(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n966), .A2(new_n969), .A3(new_n972), .ZN(G57));
endmodule


