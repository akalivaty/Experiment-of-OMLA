//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n216), .B2(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(new_n213), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT67), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(G223), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n252), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n248), .ZN(new_n257));
  INV_X1    g0057(.A(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n256), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n247), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT65), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G33), .A3(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(new_n244), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(G274), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n268), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G226), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n261), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(G179), .ZN(new_n277));
  INV_X1    g0077(.A(G1), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n213), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT68), .B1(new_n280), .B2(new_n282), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n285), .A2(new_n286), .B1(new_n278), .B2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n203), .A2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G150), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n250), .A2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n289), .B(new_n291), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n295), .A2(new_n282), .B1(new_n202), .B2(new_n280), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n276), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n277), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(G200), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n297), .B(KEYINPUT9), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n261), .A2(G190), .A3(new_n274), .A4(new_n275), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n301), .A2(new_n302), .A3(new_n306), .A4(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n300), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n253), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n256), .A2(G226), .A3(new_n248), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n246), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n265), .A2(G238), .A3(new_n270), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n269), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT13), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n247), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n269), .A2(new_n312), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n298), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n314), .A2(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n322), .A2(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n323), .A3(G169), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n322), .A2(KEYINPUT71), .A3(new_n323), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT12), .B1(new_n279), .B2(G68), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n279), .A2(KEYINPUT12), .A3(G68), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n278), .B2(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n332), .A2(new_n333), .B1(new_n283), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n290), .A2(G50), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n337), .B(new_n338), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n294), .A2(new_n259), .B1(new_n214), .B2(G68), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n282), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n342), .B2(new_n341), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n331), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n344), .B1(new_n324), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n314), .A2(new_n321), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n265), .A2(G244), .A3(new_n270), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n269), .A2(new_n356), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n257), .A2(new_n229), .B1(new_n206), .B2(new_n256), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n254), .B2(G238), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n359), .B2(new_n246), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n360), .A2(G200), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n281), .A2(new_n213), .ZN(new_n362));
  INV_X1    g0162(.A(new_n292), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n293), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n362), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n280), .A2(new_n259), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n369), .B(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n259), .B1(new_n278), .B2(G20), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n283), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n368), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n360), .B2(new_n349), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n361), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n374), .B1(new_n360), .B2(new_n298), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G179), .B2(new_n360), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n308), .A2(new_n355), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n272), .A2(G1698), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G223), .B2(G1698), .ZN(new_n382));
  AND2_X1   g0182(.A1(KEYINPUT73), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT73), .A2(G33), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT3), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n382), .B1(new_n251), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G87), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n250), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n380), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n388), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT3), .A2(G33), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT73), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n250), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT73), .A2(G33), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT75), .B(new_n390), .C1(new_n396), .C2(new_n382), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n247), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n265), .A2(G232), .A3(new_n270), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n269), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(G179), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n385), .A2(new_n251), .ZN(new_n403));
  INV_X1    g0203(.A(new_n382), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n388), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n246), .B1(new_n405), .B2(KEYINPUT75), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n400), .B1(new_n406), .B2(new_n389), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n402), .B1(new_n407), .B2(new_n298), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  INV_X1    g0209(.A(G58), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n334), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n411), .B2(new_n201), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n290), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT7), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n396), .B2(new_n214), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n385), .A2(new_n416), .A3(new_n214), .A4(new_n251), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G68), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT16), .B(new_n415), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n393), .A2(new_n249), .A3(new_n394), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n251), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n416), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n334), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n421), .B1(new_n428), .B2(new_n414), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n420), .A2(new_n429), .A3(new_n282), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n292), .A2(new_n279), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n287), .B2(new_n292), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n408), .A2(new_n409), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n409), .B1(new_n408), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT76), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n408), .A2(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n408), .A2(new_n409), .A3(new_n433), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n398), .A2(G190), .A3(new_n401), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n352), .B1(new_n398), .B2(new_n401), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n430), .A2(new_n432), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT17), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n398), .A2(G190), .A3(new_n401), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n407), .B2(new_n352), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n448), .A2(new_n433), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n436), .A2(new_n441), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n379), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT85), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n249), .B1(new_n393), .B2(new_n394), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n214), .B(G68), .C1(new_n455), .C2(new_n391), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT19), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n214), .B1(new_n316), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT82), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n387), .A2(new_n205), .A3(new_n206), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT82), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n214), .C1(new_n316), .C2(new_n457), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT19), .B1(new_n293), .B2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n282), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n366), .A2(new_n279), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT83), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  AOI211_X1 g0271(.A(new_n471), .B(new_n468), .C1(new_n466), .C2(new_n282), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n362), .B(new_n279), .C1(G1), .C2(new_n250), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n283), .B(KEYINPUT78), .C1(G1), .C2(new_n250), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n476), .A2(new_n477), .A3(G87), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(G1698), .C1(new_n455), .C2(new_n391), .ZN(new_n480));
  OAI211_X1 g0280(.A(G238), .B(new_n248), .C1(new_n455), .C2(new_n391), .ZN(new_n481));
  INV_X1    g0281(.A(G116), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n393), .B2(new_n394), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n278), .A2(G45), .ZN(new_n486));
  MUX2_X1   g0286(.A(G274), .B(G250), .S(new_n486), .Z(new_n487));
  AOI22_X1  g0287(.A1(new_n485), .A2(new_n247), .B1(new_n265), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n479), .B1(new_n488), .B2(new_n352), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n454), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(G190), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n385), .B2(new_n251), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n464), .B1(new_n492), .B2(G68), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n362), .B1(new_n493), .B2(new_n463), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n471), .B1(new_n494), .B2(new_n468), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n467), .A2(KEYINPUT83), .A3(new_n469), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n485), .A2(new_n247), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n487), .A2(new_n265), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n478), .B1(new_n500), .B2(G200), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n501), .A3(KEYINPUT85), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n490), .A2(new_n491), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n476), .A2(new_n477), .A3(new_n366), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n470), .B2(new_n472), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n504), .C1(new_n470), .C2(new_n472), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n488), .A2(G179), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n298), .B2(new_n488), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT5), .B(G41), .ZN(new_n514));
  INV_X1    g0314(.A(new_n486), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n265), .A3(G270), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n265), .A2(G274), .A3(new_n515), .A4(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n248), .B1(new_n385), .B2(new_n251), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT3), .A2(G33), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n391), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n520), .A2(G264), .B1(G303), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n403), .A2(G257), .A3(new_n248), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT86), .ZN(new_n526));
  AOI21_X1  g0326(.A(G1698), .B1(new_n385), .B2(new_n251), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G257), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n523), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n519), .B1(new_n529), .B2(new_n247), .ZN(new_n530));
  MUX2_X1   g0330(.A(new_n279), .B(new_n474), .S(G116), .Z(new_n531));
  AOI21_X1  g0331(.A(new_n362), .B1(G20), .B2(new_n482), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n214), .C1(G33), .C2(new_n205), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n532), .A2(new_n538), .A3(KEYINPUT20), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT20), .B1(new_n532), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n531), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G169), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT21), .B1(new_n530), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n519), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n403), .A2(G264), .A3(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n522), .A2(G303), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n527), .A2(new_n526), .A3(G257), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n544), .B1(new_n550), .B2(new_n246), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n532), .A2(new_n538), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT20), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n532), .A2(new_n538), .A3(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n298), .B1(new_n557), .B2(new_n531), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n551), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n543), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G190), .B(new_n544), .C1(new_n550), .C2(new_n246), .ZN(new_n561));
  INV_X1    g0361(.A(new_n541), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n530), .C2(new_n352), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n214), .A2(G87), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n522), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n483), .A2(new_n214), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n214), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(KEYINPUT22), .A2(G87), .ZN(new_n573));
  AOI211_X1 g0373(.A(G20), .B(new_n573), .C1(new_n385), .C2(new_n251), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT24), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n403), .A2(KEYINPUT22), .A3(new_n214), .A4(G87), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n483), .A2(new_n214), .B1(new_n569), .B2(new_n570), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n566), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n282), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n476), .A2(new_n477), .A3(G107), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n280), .A2(new_n206), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT25), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n403), .A2(G250), .A3(new_n248), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n395), .A2(G294), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(G1698), .C1(new_n455), .C2(new_n391), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n247), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n516), .A2(new_n265), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G264), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n518), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n325), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n592), .A2(new_n247), .B1(G264), .B2(new_n594), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n298), .B1(new_n598), .B2(new_n518), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n588), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n519), .A2(new_n325), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n541), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n549), .A2(new_n548), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n246), .B1(new_n603), .B2(new_n523), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n560), .A2(new_n563), .A3(new_n600), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT6), .B1(new_n207), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT6), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n610), .A2(new_n205), .A3(G107), .ZN(new_n611));
  OAI21_X1  g0411(.A(G20), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR4_X1   g0412(.A1(new_n259), .A2(KEYINPUT77), .A3(G20), .A4(G33), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT77), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n290), .B2(G77), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n206), .B1(new_n424), .B2(new_n427), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n282), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n476), .A2(new_n477), .A3(G97), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n280), .A2(new_n205), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n516), .A2(new_n265), .A3(G257), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n518), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(G250), .B(G1698), .C1(new_n521), .C2(new_n391), .ZN(new_n626));
  AND2_X1   g0426(.A1(KEYINPUT4), .A2(G244), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n248), .B(new_n627), .C1(new_n521), .C2(new_n391), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n628), .A3(new_n537), .ZN(new_n629));
  OAI211_X1 g0429(.A(G244), .B(new_n248), .C1(new_n455), .C2(new_n391), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT4), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n625), .B(G190), .C1(new_n632), .C2(new_n246), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT80), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n632), .B2(new_n246), .ZN(new_n635));
  INV_X1    g0435(.A(G244), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n385), .B2(new_n251), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT4), .B1(new_n637), .B2(new_n248), .ZN(new_n638));
  OAI211_X1 g0438(.A(KEYINPUT80), .B(new_n247), .C1(new_n638), .C2(new_n629), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n624), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n622), .B(new_n633), .C1(new_n640), .C2(new_n352), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n596), .A2(G200), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n586), .B1(new_n580), .B2(new_n282), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n598), .A2(G190), .A3(new_n518), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n629), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n636), .B(G1698), .C1(new_n385), .C2(new_n251), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(KEYINPUT4), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT80), .B1(new_n648), .B2(new_n247), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n632), .A2(new_n634), .A3(new_n246), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n325), .B(new_n625), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n625), .B1(new_n632), .B2(new_n246), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n298), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT81), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n422), .A2(new_n423), .B1(new_n426), .B2(new_n416), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n612), .B(new_n616), .C1(new_n656), .C2(new_n206), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n282), .B1(new_n205), .B2(new_n280), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n620), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n655), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n641), .B(new_n645), .C1(new_n654), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n607), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n453), .A2(new_n513), .A3(new_n663), .ZN(G372));
  NAND2_X1  g0464(.A1(new_n510), .A2(new_n505), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n605), .B1(new_n543), .B2(new_n559), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n600), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n479), .B1(new_n470), .B2(new_n472), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT87), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n671), .B(new_n479), .C1(new_n470), .C2(new_n472), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n500), .A2(G200), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n491), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n666), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n654), .A2(new_n622), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n677), .A3(new_n665), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n654), .A2(new_n661), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n503), .A2(new_n511), .A3(KEYINPUT26), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n453), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n434), .A2(new_n435), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n350), .A2(new_n353), .ZN(new_n687));
  INV_X1    g0487(.A(new_n378), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n348), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT17), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n449), .B1(new_n448), .B2(new_n433), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n686), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n305), .A2(new_n307), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n300), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n695), .ZN(G369));
  NAND2_X1  g0496(.A1(new_n560), .A2(new_n606), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n278), .A2(new_n214), .A3(G13), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT88), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT88), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n704), .A3(G213), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n702), .A2(new_n704), .A3(KEYINPUT89), .A4(G213), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G343), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n562), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n697), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n667), .B1(new_n562), .B2(new_n709), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n541), .B1(new_n551), .B2(G200), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n711), .A2(new_n712), .B1(new_n561), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT90), .B(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT91), .B1(new_n600), .B2(new_n709), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n596), .A2(G169), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n598), .A2(G179), .A3(new_n518), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n643), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT91), .ZN(new_n722));
  INV_X1    g0522(.A(new_n709), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n588), .A2(new_n723), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(new_n645), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n718), .A2(new_n724), .B1(new_n726), .B2(new_n600), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n718), .A2(new_n724), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n600), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n667), .A2(new_n723), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(new_n721), .B2(new_n709), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n210), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n460), .A2(G116), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(G1), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n218), .B2(new_n738), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT92), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  AND4_X1   g0543(.A1(KEYINPUT26), .A2(new_n675), .A3(new_n665), .A4(new_n677), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n503), .A2(new_n511), .A3(new_n681), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(new_n679), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n662), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n667), .A2(new_n600), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n675), .A2(new_n665), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n665), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT29), .B(new_n709), .C1(new_n746), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n723), .B1(new_n676), .B2(new_n683), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(KEYINPUT29), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n593), .A2(new_n595), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n604), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n601), .B(new_n625), .C1(new_n246), .C2(new_n632), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n488), .A4(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n625), .B1(new_n649), .B2(new_n650), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n488), .A2(G179), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n760), .A2(new_n596), .A3(new_n551), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT30), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n598), .B(new_n488), .C1(new_n550), .C2(new_n246), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n757), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n759), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n723), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT31), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n762), .A2(new_n765), .A3(KEYINPUT93), .ZN(new_n770));
  AOI21_X1  g0570(.A(KEYINPUT93), .B1(new_n762), .B2(new_n765), .ZN(new_n771));
  INV_X1    g0571(.A(new_n759), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n709), .A2(new_n768), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n769), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n512), .A2(new_n607), .A3(new_n662), .A4(new_n723), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n716), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n754), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n743), .B1(new_n780), .B2(G1), .ZN(G364));
  INV_X1    g0581(.A(G13), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n278), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n737), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n714), .B2(new_n716), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n714), .A2(new_n716), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n714), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n786), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n213), .B1(G20), .B2(new_n298), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n214), .A2(new_n325), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n349), .A3(new_n352), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n214), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n801), .A2(new_n325), .A3(new_n352), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n256), .B1(new_n259), .B2(new_n799), .C1(new_n803), .C2(new_n334), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(G190), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n214), .A2(G179), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n808), .A2(G190), .A3(G200), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n807), .A2(new_n410), .B1(new_n809), .B2(new_n387), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n808), .A2(new_n349), .A3(G200), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n206), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n805), .A2(new_n352), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n202), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n804), .A2(new_n810), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OR3_X1    g0616(.A1(KEYINPUT95), .A2(G179), .A3(G200), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT95), .B1(G179), .B2(G200), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n801), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT96), .B(G159), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n822), .A2(KEYINPUT32), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n349), .B1(new_n817), .B2(new_n818), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n214), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G97), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n822), .A2(KEYINPUT32), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n816), .A2(new_n823), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  INV_X1    g0630(.A(G303), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n811), .B1(new_n809), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G326), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n814), .A2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n832), .B(new_n834), .C1(G322), .C2(new_n806), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n826), .A2(G294), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n819), .A2(G329), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n799), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT33), .B(G317), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n256), .B(new_n839), .C1(new_n802), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n797), .B1(new_n829), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n792), .A2(new_n796), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n256), .A2(new_n210), .ZN(new_n845));
  INV_X1    g0645(.A(G355), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n845), .A2(new_n846), .B1(G116), .B2(new_n210), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT94), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n242), .A2(G45), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n403), .A2(new_n736), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(G45), .B2(new_n218), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n795), .B(new_n843), .C1(new_n844), .C2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n787), .A2(new_n789), .B1(new_n794), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NAND2_X1  g0655(.A1(new_n688), .A2(new_n709), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n361), .A2(new_n375), .B1(new_n374), .B2(new_n709), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n378), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT99), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n753), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n859), .ZN(new_n862));
  INV_X1    g0662(.A(new_n683), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n709), .B(new_n862), .C1(new_n863), .C2(new_n751), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n778), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n861), .A2(new_n778), .A3(new_n864), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n795), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n862), .A2(new_n791), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n811), .A2(new_n387), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n814), .A2(new_n831), .B1(new_n809), .B2(new_n206), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(G294), .C2(new_n806), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n819), .A2(G311), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n522), .B1(new_n799), .B2(new_n482), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G283), .B2(new_n802), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n827), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n809), .ZN(new_n878));
  INV_X1    g0678(.A(new_n811), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(G50), .B1(new_n879), .B2(G68), .ZN(new_n880));
  INV_X1    g0680(.A(new_n799), .ZN(new_n881));
  AOI22_X1  g0681(.A1(G150), .A2(new_n802), .B1(new_n881), .B2(new_n821), .ZN(new_n882));
  INV_X1    g0682(.A(G137), .ZN(new_n883));
  INV_X1    g0683(.A(G143), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n882), .B1(new_n883), .B2(new_n814), .C1(new_n884), .C2(new_n807), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT34), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n880), .B1(new_n410), .B2(new_n825), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  INV_X1    g0688(.A(new_n819), .ZN(new_n889));
  INV_X1    g0689(.A(G132), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n403), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT98), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n877), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n796), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n797), .A2(new_n791), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT97), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(G77), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n786), .B1(new_n870), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n869), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT100), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(G384));
  NOR2_X1   g0704(.A1(new_n783), .A2(new_n278), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n420), .A2(new_n282), .ZN(new_n906));
  INV_X1    g0706(.A(new_n421), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT7), .B1(new_n403), .B2(G20), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(G68), .A3(new_n418), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(new_n415), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n432), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n707), .A2(new_n708), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n452), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n398), .A2(new_n401), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(G200), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n917), .A2(new_n430), .A3(new_n432), .A4(new_n447), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n433), .A2(new_n912), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n437), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n408), .A2(new_n911), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n913), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT38), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT37), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n920), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n919), .B1(new_n451), .B2(new_n686), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n345), .A2(new_n346), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n324), .A2(G169), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n935), .A2(KEYINPUT14), .B1(new_n351), .B2(G179), .ZN(new_n936));
  INV_X1    g0736(.A(new_n330), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT71), .B1(new_n322), .B2(new_n323), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n934), .B(new_n723), .C1(new_n939), .C2(new_n354), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n345), .A2(new_n346), .A3(new_n723), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n687), .B(new_n941), .C1(new_n331), .C2(new_n347), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n859), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n766), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n769), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n777), .B2(new_n945), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n932), .A2(new_n933), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n438), .A2(new_n440), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n692), .B1(new_n949), .B2(KEYINPUT76), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n913), .B1(new_n950), .B2(new_n441), .ZN(new_n951));
  INV_X1    g0751(.A(new_n925), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n927), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n946), .B1(new_n926), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n948), .B1(new_n954), .B2(KEYINPUT40), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n769), .A2(new_n944), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n663), .A2(new_n513), .A3(new_n709), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI221_X4 g0758(.A(new_n927), .B1(new_n921), .B2(new_n924), .C1(new_n452), .C2(new_n914), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT38), .B1(new_n915), .B2(new_n925), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n943), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(KEYINPUT103), .A3(new_n933), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n947), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT104), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n453), .A2(new_n958), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n715), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n964), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT101), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n953), .A2(new_n926), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n940), .A2(new_n942), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n723), .B(new_n859), .C1(new_n676), .C2(new_n683), .ZN(new_n972));
  INV_X1    g0772(.A(new_n856), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n970), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n686), .A2(new_n912), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n969), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n926), .A2(new_n931), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT39), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n953), .A2(KEYINPUT39), .A3(new_n926), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n348), .A2(new_n709), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT102), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n974), .A2(new_n969), .A3(new_n976), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n752), .B(new_n453), .C1(KEYINPUT29), .C2(new_n753), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n695), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n905), .B1(new_n968), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n992), .B2(new_n968), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n609), .A2(new_n611), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n482), .B(new_n216), .C1(new_n996), .C2(KEYINPUT35), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(KEYINPUT35), .B2(new_n996), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT36), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n218), .A2(new_n259), .A3(new_n411), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n334), .A2(G50), .ZN(new_n1001));
  OAI211_X1 g0801(.A(G1), .B(new_n782), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n994), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT105), .ZN(G367));
  INV_X1    g0804(.A(new_n850), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n844), .B1(new_n210), .B2(new_n365), .C1(new_n1005), .C2(new_n235), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(new_n786), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n709), .B1(new_n670), .B2(new_n672), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n666), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n750), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n811), .A2(new_n259), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n814), .A2(new_n884), .B1(new_n809), .B2(new_n410), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G150), .C2(new_n806), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n256), .B1(new_n799), .B2(new_n202), .C1(new_n803), .C2(new_n820), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G137), .B2(new_n819), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(new_n334), .C2(new_n825), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n799), .A2(new_n830), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n403), .B(new_n1017), .C1(G294), .C2(new_n802), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n809), .A2(new_n482), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G317), .A2(new_n819), .B1(new_n1019), .B2(KEYINPUT46), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(KEYINPUT46), .C2(new_n1019), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n811), .A2(new_n205), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G303), .B2(new_n806), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n838), .B2(new_n814), .C1(new_n206), .C2(new_n825), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1016), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n1007), .B1(new_n1010), .B2(new_n793), .C1(new_n1026), .C2(new_n797), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT109), .Z(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n658), .A2(new_n620), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n723), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n654), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n651), .B(new_n653), .C1(new_n659), .C2(new_n660), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n641), .A3(new_n1031), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT106), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT106), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1036), .A3(new_n641), .A4(new_n1031), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1032), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n734), .A2(new_n1039), .A3(KEYINPUT45), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT45), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n733), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n727), .A2(new_n1042), .B1(new_n600), .B2(new_n723), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1043), .B2(new_n1038), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n734), .B2(new_n1039), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1043), .A2(new_n1038), .A3(new_n1046), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n728), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1052), .A2(new_n729), .A3(new_n1049), .A4(new_n1048), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n732), .A2(new_n733), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n727), .A2(new_n1042), .ZN(new_n1057));
  AND4_X1   g0857(.A1(new_n716), .A2(new_n1056), .A3(new_n714), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1056), .A2(new_n1057), .B1(new_n714), .B2(new_n716), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n754), .A2(new_n1060), .A3(new_n778), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT108), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT108), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1054), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n780), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n737), .B(KEYINPUT41), .Z(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n785), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1056), .A2(new_n1038), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT42), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1033), .B1(new_n1038), .B2(new_n600), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n709), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1071), .A2(new_n1073), .B1(KEYINPUT43), .B2(new_n1010), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n728), .A2(new_n1039), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1029), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT110), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1079), .B(new_n1080), .ZN(G387));
  NAND2_X1  g0881(.A1(new_n1061), .A2(new_n737), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT113), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT113), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1061), .A2(new_n1084), .A3(new_n737), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(new_n780), .C2(new_n1060), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n727), .A2(new_n792), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n845), .A2(new_n739), .B1(G107), .B2(new_n210), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n232), .A2(new_n267), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n739), .ZN(new_n1090));
  AOI211_X1 g0890(.A(G45), .B(new_n1090), .C1(G68), .C2(G77), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n292), .A2(G50), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT50), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1005), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1088), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n844), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n786), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(G159), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n202), .A2(new_n807), .B1(new_n814), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1022), .B(new_n1099), .C1(G77), .C2(new_n878), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n826), .A2(new_n366), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT111), .B(G150), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n819), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n799), .A2(new_n334), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n396), .B(new_n1104), .C1(new_n363), .C2(new_n802), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n403), .B1(G116), .B2(new_n879), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G311), .A2(new_n802), .B1(new_n881), .B2(G303), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n806), .A2(G317), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT112), .B(G322), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n1109), .C1(new_n814), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT48), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n826), .A2(G283), .B1(G294), .B2(new_n878), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT49), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1107), .B1(new_n833), .B2(new_n889), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1106), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1097), .B1(new_n1120), .B2(new_n796), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1060), .A2(new_n785), .B1(new_n1087), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1086), .A2(new_n1122), .ZN(G393));
  NAND3_X1  g0923(.A1(new_n1051), .A2(KEYINPUT114), .A3(new_n1053), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT114), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1125), .B(new_n728), .C1(new_n1045), .C2(new_n1050), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n737), .B1(new_n1062), .B2(new_n1127), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n844), .B1(new_n205), .B2(new_n210), .C1(new_n1005), .C2(new_n239), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n786), .ZN(new_n1130));
  INV_X1    g0930(.A(G294), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n522), .B1(new_n1131), .B2(new_n799), .C1(new_n803), .C2(new_n831), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n812), .B(new_n1132), .C1(G283), .C2(new_n878), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n806), .A2(G311), .B1(new_n813), .B2(G317), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT52), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n826), .A2(G116), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n889), .A2(new_n1110), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n806), .A2(G159), .B1(new_n813), .B2(G150), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT51), .Z(new_n1140));
  INV_X1    g0940(.A(new_n871), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n826), .A2(G77), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n799), .A2(new_n292), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n396), .B(new_n1143), .C1(G50), .C2(new_n802), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n819), .A2(G143), .B1(new_n878), .B2(G68), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT116), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1138), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1130), .B1(new_n1148), .B2(new_n796), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1039), .B2(new_n793), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n784), .B1(new_n1127), .B2(KEYINPUT115), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT115), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1124), .A2(new_n1153), .A3(new_n1126), .ZN(new_n1154));
  AOI211_X1 g0954(.A(KEYINPUT117), .B(new_n1151), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT117), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1127), .A2(KEYINPUT115), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n785), .A3(new_n1154), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1158), .B2(new_n1150), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1128), .B1(new_n1155), .B2(new_n1159), .ZN(G390));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n256), .B1(new_n799), .B2(new_n1161), .C1(new_n803), .C2(new_n883), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n878), .A2(new_n1102), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G125), .C2(new_n819), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n813), .A2(G128), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n202), .B2(new_n811), .C1(new_n807), .C2(new_n890), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G159), .B2(new_n826), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n522), .B1(new_n205), .B2(new_n799), .C1(new_n803), .C2(new_n206), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n482), .A2(new_n807), .B1(new_n814), .B2(new_n830), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n334), .A2(new_n811), .B1(new_n809), .B2(new_n387), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n889), .A2(new_n1131), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1165), .A2(new_n1168), .B1(new_n1142), .B2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n786), .B1(new_n363), .B2(new_n899), .C1(new_n1174), .C2(new_n797), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n982), .B2(new_n790), .ZN(new_n1176));
  INV_X1    g0976(.A(G330), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n956), .B2(new_n957), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n943), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n971), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n864), .B2(new_n856), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n984), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n982), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n858), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n745), .A2(new_n679), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT26), .A4(new_n665), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n723), .B(new_n1184), .C1(new_n676), .C2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n971), .B1(new_n1188), .B2(new_n973), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n978), .A2(new_n984), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1179), .B1(new_n1183), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT118), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(new_n984), .B1(new_n980), .B2(new_n981), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n716), .B(new_n943), .C1(new_n776), .C2(new_n777), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n709), .B(new_n858), .C1(new_n746), .C2(new_n751), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1180), .B1(new_n1198), .B2(new_n856), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1199), .B2(new_n1190), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1197), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(KEYINPUT118), .A3(new_n1183), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1193), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1176), .B1(new_n1205), .B2(new_n785), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n453), .A2(new_n1178), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n990), .A2(new_n695), .A3(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n716), .B(new_n862), .C1(new_n776), .C2(new_n777), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1209), .A2(new_n1180), .B1(new_n1178), .B2(new_n943), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n972), .A2(new_n973), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1198), .A2(new_n1197), .A3(new_n856), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n971), .B1(new_n1178), .B2(new_n860), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1208), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n737), .B1(new_n1205), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1183), .A2(new_n1192), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1179), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1196), .A2(new_n1200), .A3(new_n1194), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT118), .B1(new_n1203), .B2(new_n1183), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1216), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(KEYINPUT119), .B(new_n1206), .C1(new_n1217), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n990), .A2(new_n695), .A3(new_n1207), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1210), .A2(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n737), .A3(new_n1223), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT119), .B1(new_n1232), .B2(new_n1206), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1226), .A2(new_n1233), .ZN(G378));
  INV_X1    g1034(.A(new_n947), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n946), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n948), .B(KEYINPUT40), .C1(new_n970), .C2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT103), .B1(new_n961), .B2(new_n933), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G330), .B(new_n1235), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1240));
  XNOR2_X1  g1040(.A(new_n308), .B(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n912), .A2(new_n297), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT122), .Z(new_n1243));
  XOR2_X1   g1043(.A(new_n1241), .B(new_n1243), .Z(new_n1244));
  NOR2_X1   g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1244), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n963), .B2(G330), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n989), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n987), .A2(new_n977), .A3(new_n985), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n963), .A2(G330), .A3(new_n1246), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1248), .A2(new_n1252), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT123), .B1(new_n1253), .B2(KEYINPUT57), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n738), .B1(new_n1253), .B2(KEYINPUT57), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1250), .A2(new_n1251), .B1(new_n988), .B2(new_n986), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1208), .B1(new_n1205), .B2(new_n1216), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1256), .B(new_n1257), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1254), .A2(new_n1255), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1244), .A2(new_n790), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n786), .B1(new_n899), .B2(G50), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n403), .A2(G41), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(G33), .A2(G41), .ZN(new_n1267));
  OR3_X1    g1067(.A1(new_n1266), .A2(G50), .A3(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G97), .A2(new_n802), .B1(new_n881), .B2(new_n366), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1269), .B(new_n1266), .C1(new_n259), .C2(new_n809), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n806), .A2(G107), .B1(new_n813), .B2(G116), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n410), .B2(new_n811), .C1(new_n334), .C2(new_n825), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1270), .B(new_n1272), .C1(G283), .C2(new_n819), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1268), .B1(new_n1273), .B2(KEYINPUT58), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT120), .Z(new_n1275));
  AND2_X1   g1075(.A1(new_n813), .A2(G125), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n803), .A2(new_n890), .B1(new_n883), .B2(new_n799), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(G128), .C2(new_n806), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n809), .A2(new_n1161), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT121), .ZN(new_n1280));
  INV_X1    g1080(.A(G150), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1278), .B(new_n1280), .C1(new_n1281), .C2(new_n825), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(KEYINPUT59), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n819), .A2(G124), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1284), .B(new_n1267), .C1(new_n811), .C2(new_n820), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n1282), .B2(KEYINPUT59), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1283), .A2(new_n1286), .B1(KEYINPUT58), .B2(new_n1273), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1275), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1265), .B1(new_n1288), .B2(new_n796), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1264), .A2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1260), .B2(new_n784), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1263), .A2(new_n1292), .ZN(G375));
  INV_X1    g1093(.A(new_n1229), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1208), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1068), .A3(new_n1230), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1229), .A2(KEYINPUT124), .A3(new_n785), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n786), .B1(new_n899), .B2(G68), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1101), .B1(new_n830), .B2(new_n807), .ZN(new_n1299));
  XOR2_X1   g1099(.A(new_n1299), .B(KEYINPUT125), .Z(new_n1300));
  OAI221_X1 g1100(.A(new_n522), .B1(new_n206), .B2(new_n799), .C1(new_n803), .C2(new_n482), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1011), .B1(G294), .B2(new_n813), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n205), .B2(new_n809), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1301), .B(new_n1303), .C1(G303), .C2(new_n819), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n825), .A2(new_n202), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n890), .A2(new_n814), .B1(new_n807), .B2(new_n883), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n410), .A2(new_n811), .B1(new_n809), .B2(new_n1098), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n819), .A2(G128), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n803), .A2(new_n1161), .B1(new_n1281), .B2(new_n799), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(new_n396), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1309), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1305), .B1(new_n1306), .B2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1298), .B1(new_n1314), .B2(new_n796), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n971), .B2(new_n791), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1294), .B2(new_n784), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1296), .A2(new_n1297), .A3(new_n1316), .A4(new_n1318), .ZN(G381));
  AND3_X1   g1119(.A1(new_n1086), .A2(new_n854), .A3(new_n1122), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OR3_X1    g1121(.A1(new_n1321), .A2(G384), .A3(G381), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1232), .A2(new_n1206), .ZN(new_n1323));
  OR3_X1    g1123(.A1(new_n1322), .A2(G390), .A3(new_n1323), .ZN(new_n1324));
  OR3_X1    g1124(.A1(new_n1324), .A2(G387), .A3(G375), .ZN(G407));
  INV_X1    g1125(.A(new_n1323), .ZN(new_n1326));
  INV_X1    g1126(.A(G213), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1327), .A2(G343), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G407), .B(G213), .C1(G375), .C2(new_n1329), .ZN(G409));
  NAND3_X1  g1130(.A1(new_n1263), .A2(G378), .A3(new_n1292), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1260), .A2(new_n1067), .A3(new_n1261), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1326), .B1(new_n1332), .B2(new_n1291), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1328), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1318), .A2(new_n1297), .A3(new_n1316), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1212), .A2(new_n1215), .A3(KEYINPUT60), .A4(new_n1208), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n737), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1230), .A2(KEYINPUT60), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1295), .B2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(G384), .B1(new_n1336), .B2(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1336), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n902), .B(KEYINPUT100), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1334), .A2(new_n1335), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(KEYINPUT62), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1328), .A2(G2897), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1345), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1349), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1341), .A2(new_n1344), .A3(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1348), .A2(new_n1350), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1328), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT62), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(new_n1356), .A3(new_n1345), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1347), .A2(new_n1353), .A3(new_n1354), .A4(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n854), .B1(new_n1086), .B2(new_n1122), .ZN(new_n1359));
  OR2_X1    g1159(.A1(new_n1320), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G390), .A2(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1080), .B1(new_n1320), .B2(new_n1359), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1362), .B(new_n1128), .C1(new_n1155), .C2(new_n1159), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1361), .A2(new_n1079), .A3(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1079), .B1(new_n1361), .B2(new_n1363), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1358), .A2(new_n1367), .ZN(new_n1368));
  NOR3_X1   g1168(.A1(new_n1364), .A2(new_n1365), .A3(KEYINPUT61), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT126), .ZN(new_n1370));
  AND3_X1   g1170(.A1(new_n1341), .A2(new_n1344), .A3(new_n1351), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1351), .B1(new_n1341), .B2(new_n1344), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1370), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1350), .A2(KEYINPUT126), .A3(new_n1352), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1369), .B1(new_n1355), .B2(new_n1375), .ZN(new_n1376));
  AOI21_X1  g1176(.A(KEYINPUT63), .B1(new_n1355), .B2(new_n1345), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1355), .A2(KEYINPUT63), .A3(new_n1345), .ZN(new_n1379));
  AOI21_X1  g1179(.A(KEYINPUT127), .B1(new_n1378), .B2(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1361), .A2(new_n1363), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1079), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1361), .A2(new_n1363), .A3(new_n1079), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1383), .A2(new_n1354), .A3(new_n1384), .ZN(new_n1385));
  AND2_X1   g1185(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1386));
  AOI21_X1  g1186(.A(new_n1385), .B1(new_n1348), .B2(new_n1386), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT63), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1346), .A2(new_n1388), .ZN(new_n1389));
  AND4_X1   g1189(.A1(KEYINPUT127), .A2(new_n1387), .A3(new_n1379), .A4(new_n1389), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1368), .B1(new_n1380), .B2(new_n1390), .ZN(G405));
  NAND2_X1  g1191(.A1(G375), .A2(new_n1326), .ZN(new_n1392));
  AND2_X1   g1192(.A1(new_n1392), .A2(new_n1331), .ZN(new_n1393));
  OR2_X1    g1193(.A1(new_n1393), .A2(new_n1345), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1393), .A2(new_n1345), .ZN(new_n1395));
  AND3_X1   g1195(.A1(new_n1394), .A2(new_n1395), .A3(new_n1366), .ZN(new_n1396));
  AOI21_X1  g1196(.A(new_n1366), .B1(new_n1394), .B2(new_n1395), .ZN(new_n1397));
  NOR2_X1   g1197(.A1(new_n1396), .A2(new_n1397), .ZN(G402));
endmodule


