//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203));
  AOI21_X1  g002(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT72), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n203), .B1(new_n208), .B2(KEYINPUT73), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n210), .A3(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n206), .A2(new_n210), .A3(new_n203), .A4(new_n207), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n212), .B2(new_n214), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT76), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n220), .A2(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n219), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  AND4_X1   g035(.A1(KEYINPUT25), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(new_n221), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n226), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT65), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT25), .A4(new_n234), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n221), .B1(new_n225), .B2(new_n227), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n236), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT27), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G183gat), .ZN(new_n251));
  INV_X1    g050(.A(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT27), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n249), .B1(new_n252), .B2(KEYINPUT27), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n248), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT28), .A4(new_n256), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n229), .A2(new_n230), .ZN(new_n261));
  INV_X1    g060(.A(new_n234), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(KEYINPUT26), .ZN(new_n263));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT26), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n267), .A2(new_n224), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT29), .B1(new_n247), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT75), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n218), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n262), .B1(KEYINPUT23), .B2(new_n264), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n219), .B1(new_n261), .B2(new_n232), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n241), .A2(KEYINPUT65), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n245), .B1(new_n243), .B2(new_n244), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n279), .A2(new_n236), .B1(new_n260), .B2(new_n268), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT76), .B(new_n274), .C1(new_n280), .C2(KEYINPUT29), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n247), .A2(new_n269), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g085(.A(KEYINPUT77), .B(new_n271), .C1(new_n247), .C2(new_n269), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n217), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT78), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT77), .B1(new_n280), .B2(new_n271), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n223), .A2(new_n220), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n225), .A2(new_n227), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n235), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n277), .A2(new_n278), .B1(new_n296), .B2(new_n219), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n267), .A2(new_n224), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n258), .B2(new_n259), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n283), .B(new_n285), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n281), .A3(new_n273), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n217), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(new_n304), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n270), .A2(KEYINPUT79), .A3(new_n285), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n212), .A2(new_n214), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT79), .B1(new_n270), .B2(new_n285), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n284), .A2(new_n272), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n306), .A2(new_n308), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n305), .A2(KEYINPUT30), .A3(new_n311), .A4(new_n315), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n302), .A2(new_n303), .A3(new_n217), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n303), .B1(new_n302), .B2(new_n217), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n314), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT0), .ZN(new_n324));
  XNOR2_X1  g123(.A(G57gat), .B(G85gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333));
  NAND2_X1  g132(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n332), .A2(new_n333), .A3(G120gat), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G113gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n333), .B1(new_n341), .B2(G120gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n331), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G113gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n328), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G155gat), .B(G162gat), .ZN(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  INV_X1    g152(.A(G162gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT2), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  INV_X1    g156(.A(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n343), .A2(new_n348), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n332), .A2(G120gat), .A3(new_n334), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n337), .A3(new_n335), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n347), .B1(new_n372), .B2(new_n331), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT84), .B1(new_n373), .B2(new_n367), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n366), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n335), .A2(new_n337), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n330), .B1(new_n377), .B2(new_n371), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n375), .B(new_n376), .C1(new_n378), .C2(new_n347), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n369), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n381), .B(KEYINPUT82), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT5), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT81), .B(new_n387), .C1(new_n356), .C2(new_n366), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n343), .A2(new_n348), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n382), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n368), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n397), .A3(KEYINPUT83), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT81), .B1(new_n367), .B2(new_n387), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n376), .A2(new_n385), .A3(KEYINPUT3), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n367), .A2(new_n387), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n399), .A2(new_n391), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(new_n394), .A3(new_n395), .A4(new_n383), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n384), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(KEYINPUT85), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(new_n395), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n382), .A2(KEYINPUT5), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n407), .A2(new_n402), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n327), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n374), .A2(new_n379), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n368), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n416), .B2(new_n382), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT83), .B1(new_n392), .B2(new_n397), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n404), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n326), .A3(new_n411), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n413), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT6), .B(new_n327), .C1(new_n406), .C2(new_n412), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n311), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n423), .A2(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n322), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n321), .B1(new_n316), .B2(new_n320), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n202), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n316), .A2(new_n320), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n432), .A2(KEYINPUT86), .A3(new_n322), .A4(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(G228gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n401), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n307), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT87), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n212), .A2(new_n214), .A3(new_n439), .A4(new_n435), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n438), .A2(new_n387), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n434), .B(new_n437), .C1(new_n441), .C2(new_n367), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n308), .A2(new_n435), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n367), .B1(new_n443), .B2(new_n387), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n436), .B1(new_n215), .B2(new_n216), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT88), .B(new_n436), .C1(new_n215), .C2(new_n216), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n442), .B1(new_n449), .B2(new_n434), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT31), .B(G50gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(G22gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n442), .B(new_n454), .C1(new_n449), .C2(new_n434), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT69), .B(new_n391), .C1(new_n297), .C2(new_n299), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n280), .B2(new_n373), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n280), .A2(new_n373), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT33), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(KEYINPUT32), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n464), .B2(new_n466), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT70), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n471), .ZN(new_n477));
  INV_X1    g276(.A(new_n470), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n467), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n473), .A2(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n465), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n483), .B(KEYINPUT34), .Z(new_n484));
  OR2_X1    g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n481), .ZN(new_n486));
  INV_X1    g285(.A(new_n477), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n476), .B1(new_n475), .B2(new_n471), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n486), .B(new_n484), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n459), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n430), .A2(new_n433), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT35), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n423), .A2(new_n424), .ZN(new_n494));
  AND4_X1   g293(.A1(new_n493), .A2(new_n494), .A3(new_n457), .A4(new_n456), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n482), .A2(new_n484), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n498), .A3(new_n484), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n425), .A2(new_n426), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n316), .A3(new_n320), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n495), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n492), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n497), .A2(new_n499), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n485), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n485), .A2(KEYINPUT36), .A3(new_n489), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(new_n311), .C1(new_n317), .C2(new_n318), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n302), .A2(new_n217), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n307), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n513), .B(new_n314), .C1(new_n512), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT38), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n319), .B2(KEYINPUT37), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(new_n314), .A3(new_n513), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n407), .A2(new_n402), .A3(new_n409), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n382), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT39), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n380), .B2(new_n383), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n327), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n528), .A3(new_n382), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT40), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n413), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT40), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n458), .B1(new_n502), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n510), .A2(new_n511), .B1(new_n525), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n430), .A2(new_n433), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n458), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n506), .A2(new_n540), .A3(KEYINPUT89), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT89), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n511), .B1(new_n500), .B2(KEYINPUT36), .ZN(new_n543));
  INV_X1    g342(.A(new_n536), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n523), .B1(new_n519), .B2(new_n521), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n459), .B1(new_n430), .B2(new_n433), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n504), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n542), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G1gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554));
  MUX2_X1   g353(.A(G1gat), .B(new_n553), .S(new_n554), .Z(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(G8gat), .Z(new_n556));
  XOR2_X1   g355(.A(G57gat), .B(G64gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  AND2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT94), .ZN(new_n563));
  INV_X1    g362(.A(new_n561), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n557), .C1(KEYINPUT9), .C2(new_n559), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT95), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n556), .B1(new_n567), .B2(KEYINPUT21), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n566), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT96), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT97), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n574), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(new_n577), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n570), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT98), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n575), .A2(new_n578), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n569), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n585), .B1(new_n583), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n568), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(new_n568), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n592), .B2(new_n595), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(KEYINPUT91), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(KEYINPUT91), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(G29gat), .A2(G36gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G50gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G43gat), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(G43gat), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n607), .A2(KEYINPUT15), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n609), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT15), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n614), .ZN(new_n616));
  INV_X1    g415(.A(new_n602), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n603), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n615), .A2(new_n616), .A3(new_n606), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT17), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G85gat), .A2(G92gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(KEYINPUT101), .A3(KEYINPUT7), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(KEYINPUT7), .B2(new_n626), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT101), .B1(new_n626), .B2(KEYINPUT7), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G99gat), .B(G106gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n634), .A2(new_n620), .B1(KEYINPUT41), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n641), .A2(new_n643), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT100), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n601), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G230gat), .ZN(new_n654));
  INV_X1    g453(.A(G233gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n634), .A2(new_n563), .A3(new_n565), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n567), .B2(new_n634), .ZN(new_n658));
  NOR2_X1   g457(.A1(KEYINPUT102), .A2(KEYINPUT10), .ZN(new_n659));
  AND2_X1   g458(.A1(KEYINPUT102), .A2(KEYINPUT10), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n634), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n656), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n656), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n664), .A2(new_n665), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n556), .A2(new_n620), .ZN(new_n674));
  INV_X1    g473(.A(new_n556), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n621), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(G229gat), .A2(G233gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(KEYINPUT18), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n556), .B(new_n620), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n677), .B(KEYINPUT13), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n677), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT18), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G113gat), .B(G141gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(G169gat), .B(G197gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT12), .Z(new_n693));
  OAI211_X1 g492(.A(new_n687), .B(new_n693), .C1(KEYINPUT93), .C2(new_n682), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT93), .ZN(new_n695));
  INV_X1    g494(.A(new_n693), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n683), .B(new_n686), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n673), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n551), .A2(new_n653), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n494), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n502), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n552), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n706), .A2(G8gat), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G8gat), .B1(new_n706), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n707), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n701), .B2(new_n543), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n508), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n701), .B2(new_n715), .ZN(G1326gat));
  NAND2_X1  g515(.A1(new_n702), .A2(new_n458), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT104), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT105), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n718), .B(new_n720), .ZN(G1327gat));
  NAND3_X1  g520(.A1(new_n541), .A2(new_n550), .A3(new_n652), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n601), .A2(new_n700), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(G29gat), .A3(new_n494), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT45), .Z(new_n727));
  OAI21_X1  g526(.A(new_n537), .B1(new_n539), .B2(KEYINPUT107), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n547), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n506), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n652), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n722), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT106), .B1(new_n722), .B2(KEYINPUT44), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n724), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n494), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n738), .ZN(G1328gat));
  OR2_X1    g538(.A1(new_n503), .A2(G36gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT46), .B1(new_n725), .B2(new_n740), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G36gat), .B1(new_n737), .B2(new_n503), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1329gat));
  OAI21_X1  g547(.A(G43gat), .B1(new_n737), .B2(new_n543), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n725), .A2(G43gat), .A3(new_n508), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT47), .B1(new_n751), .B2(KEYINPUT110), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n753), .B(new_n754), .C1(new_n749), .C2(new_n750), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(G1330gat));
  INV_X1    g555(.A(new_n725), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(KEYINPUT111), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n458), .B1(new_n757), .B2(KEYINPUT111), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n608), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n736), .A2(G50gat), .A3(new_n458), .A4(new_n724), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g562(.A1(new_n653), .A2(new_n699), .A3(new_n673), .A4(new_n731), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n703), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT112), .B(G57gat), .Z(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1332gat));
  AOI21_X1  g566(.A(new_n503), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n769), .B(new_n770), .Z(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n764), .A2(new_n772), .A3(new_n500), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n764), .A2(new_n510), .A3(new_n511), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n772), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g575(.A1(new_n764), .A2(new_n458), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n599), .A2(new_n600), .A3(new_n698), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n673), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n736), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(new_n494), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G85gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n782), .A2(new_n779), .A3(new_n494), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n780), .A2(new_n731), .A3(new_n652), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n780), .A2(new_n731), .A3(new_n788), .A4(new_n652), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n673), .A2(new_n623), .A3(new_n703), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n784), .A2(new_n785), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n736), .A2(new_n502), .A3(new_n781), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n624), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n673), .A2(new_n624), .A3(new_n502), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT114), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n786), .A2(new_n802), .A3(new_n788), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n786), .B1(new_n802), .B2(new_n788), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n800), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n794), .B2(G92gat), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n797), .A2(new_n801), .B1(new_n798), .B2(new_n807), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n782), .B2(new_n543), .ZN(new_n809));
  INV_X1    g608(.A(new_n673), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n810), .A2(G99gat), .A3(new_n508), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n791), .B2(new_n811), .ZN(G1338gat));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n736), .A2(new_n458), .A3(new_n781), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n810), .A2(G106gat), .A3(new_n459), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n787), .A2(new_n789), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n813), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT118), .B(new_n819), .C1(new_n814), .C2(G106gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n816), .B1(new_n803), .B2(new_n804), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n815), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(KEYINPUT53), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT117), .B(new_n818), .C1(new_n815), .C2(new_n825), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n592), .A2(new_n595), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n596), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n661), .A2(new_n662), .A3(new_n656), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n832), .A2(new_n663), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n671), .B1(new_n663), .B2(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  INV_X1    g637(.A(new_n836), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n834), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n837), .A2(new_n840), .A3(new_n698), .A4(new_n672), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n676), .A2(new_n677), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n679), .A2(new_n680), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n692), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n683), .A2(new_n696), .A3(new_n686), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n673), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n652), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n837), .A2(new_n672), .A3(new_n840), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n844), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n651), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n598), .B(new_n831), .C1(new_n847), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n673), .A2(new_n698), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n651), .B(new_n852), .C1(new_n599), .C2(new_n600), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n502), .A2(new_n494), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n508), .A2(new_n458), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n699), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n856), .A2(new_n490), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n698), .A2(new_n341), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT119), .Z(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1340gat));
  AOI21_X1  g664(.A(new_n336), .B1(new_n858), .B2(new_n673), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT120), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n861), .A2(new_n336), .A3(new_n673), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n859), .B2(new_n601), .ZN(new_n870));
  INV_X1    g669(.A(G127gat), .ZN(new_n871));
  INV_X1    g670(.A(new_n601), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n861), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n651), .A2(G134gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n856), .A2(new_n490), .A3(new_n875), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT56), .Z(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n859), .B2(new_n651), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1343gat));
  AOI21_X1  g678(.A(new_n459), .B1(new_n851), .B2(new_n853), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n543), .A2(new_n855), .ZN(new_n885));
  AND2_X1   g684(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n887), .A3(new_n698), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n884), .A2(new_n887), .A3(new_n890), .A4(new_n698), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n357), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n885), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n880), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n699), .A2(G141gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n888), .A2(G141gat), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n892), .A2(new_n898), .B1(new_n897), .B2(new_n899), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n358), .A3(new_n673), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n810), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(KEYINPUT59), .A3(new_n358), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n810), .B1(new_n881), .B2(new_n883), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n893), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n902), .B1(new_n905), .B2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n903), .B2(new_n601), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n353), .A3(new_n872), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n903), .B2(new_n651), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n894), .A2(new_n354), .A3(new_n652), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n503), .A2(new_n703), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n854), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n490), .ZN(new_n919));
  AOI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n698), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n857), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(new_n229), .A3(new_n699), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n922), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n230), .A3(new_n673), .ZN(new_n924));
  OAI21_X1  g723(.A(G176gat), .B1(new_n921), .B2(new_n810), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND4_X1  g725(.A1(new_n919), .A2(new_n251), .A3(new_n253), .A4(new_n872), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n921), .A2(new_n601), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n252), .ZN(new_n929));
  XOR2_X1   g728(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n919), .A2(new_n256), .A3(new_n652), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n918), .A2(new_n652), .A3(new_n857), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(G190gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n933), .B2(G190gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1351gat));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(G197gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n881), .A2(new_n883), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n543), .A2(new_n917), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n940), .B1(new_n943), .B2(new_n698), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n880), .A2(new_n942), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(new_n698), .A3(new_n940), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n944), .A2(new_n946), .ZN(G1352gat));
  INV_X1    g746(.A(G204gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n948), .A3(new_n673), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT62), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n907), .A2(new_n942), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n948), .ZN(G1353gat));
  INV_X1    g752(.A(G211gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n945), .A2(new_n954), .A3(new_n872), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n943), .A2(new_n872), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n943), .A2(G218gat), .A3(new_n652), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n945), .A2(new_n652), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n961), .A2(new_n962), .A3(G218gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n961), .B2(G218gat), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(G1355gat));
endmodule


