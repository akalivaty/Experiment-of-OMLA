//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT81), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n198));
  OAI21_X1  g012(.A(G128), .B1(new_n198), .B2(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(G143), .B2(new_n192), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n196), .A2(new_n200), .A3(G128), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT10), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G104), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT3), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n211), .A3(KEYINPUT3), .A4(G104), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n213), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT78), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n211), .A3(G104), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n218), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT78), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n213), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n211), .A2(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n215), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n209), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n225), .B2(new_n213), .ZN(new_n232));
  AOI211_X1 g046(.A(KEYINPUT78), .B(new_n212), .C1(new_n224), .C2(new_n218), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n209), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n208), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT64), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G134), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(G137), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(G137), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT64), .B(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n241), .B2(new_n243), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n238), .A2(new_n240), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT11), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n201), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n205), .B1(new_n259), .B2(new_n196), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n228), .A2(new_n230), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n207), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n229), .B1(new_n224), .B2(new_n218), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT0), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n196), .B1(new_n266), .B2(new_n258), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT0), .B(G128), .Z(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(new_n196), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n232), .A2(new_n233), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT4), .B1(new_n263), .B2(new_n210), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n265), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n236), .A2(new_n257), .A3(new_n262), .A4(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G110), .B(G140), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G227), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT79), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n206), .A3(new_n234), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n261), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT12), .A3(new_n256), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n256), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n279), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n236), .A2(new_n262), .A3(new_n272), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n256), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n278), .B1(new_n290), .B2(new_n273), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n190), .B(new_n191), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT12), .B1(new_n283), .B2(new_n256), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n286), .B(new_n257), .C1(new_n282), .C2(new_n261), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n273), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n277), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n273), .A2(new_n278), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n290), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(G469), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n190), .A2(new_n191), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n292), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G221), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT9), .B(G234), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n305), .B2(new_n191), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n302), .A2(KEYINPUT80), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT80), .B1(new_n302), .B2(new_n307), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G116), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G119), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT5), .ZN(new_n316));
  OAI21_X1  g130(.A(G113), .B1(new_n313), .B2(KEYINPUT5), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT2), .B(G113), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n315), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n316), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n231), .B2(new_n235), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(KEYINPUT67), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT2), .B(G113), .Z(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n318), .A3(KEYINPUT67), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n328), .B(new_n265), .C1(new_n270), .C2(new_n271), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(KEYINPUT82), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n320), .B1(new_n281), .B2(new_n234), .ZN(new_n332));
  INV_X1    g146(.A(new_n271), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n264), .B(new_n327), .C1(new_n228), .C2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G122), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n332), .A2(new_n334), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n336), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n330), .A2(new_n335), .A3(new_n340), .A4(new_n337), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n339), .B1(new_n338), .B2(new_n342), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n269), .A2(G125), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n206), .B2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G224), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT84), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n338), .A2(new_n342), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT83), .A3(new_n344), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n357));
  INV_X1    g171(.A(new_n351), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT7), .B1(new_n349), .B2(G953), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n348), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n348), .A2(new_n362), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT87), .Z(new_n365));
  AOI211_X1 g179(.A(new_n363), .B(new_n365), .C1(new_n341), .C2(new_n336), .ZN(new_n366));
  INV_X1    g180(.A(new_n280), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n367), .B(new_n320), .C1(KEYINPUT79), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n336), .B(KEYINPUT8), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT85), .B1(new_n281), .B2(new_n234), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n320), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT86), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n311), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n357), .B1(new_n356), .B2(new_n358), .ZN(new_n376));
  AOI211_X1 g190(.A(KEYINPUT84), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n311), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n189), .B(new_n310), .C1(new_n375), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n246), .B1(new_n245), .B2(new_n249), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n251), .A2(new_n254), .A3(G131), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n269), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n204), .A2(new_n205), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n248), .A2(G137), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n253), .A2(G134), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n250), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n389), .A3(KEYINPUT30), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT65), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n256), .A2(new_n393), .A3(new_n269), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n328), .B(new_n390), .C1(new_n395), .C2(KEYINPUT30), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G101), .ZN(new_n397));
  NOR2_X1   g211(.A1(G237), .A2(G953), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G210), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n384), .A2(new_n389), .A3(new_n327), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n396), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT28), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n404), .B(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n395), .A2(new_n327), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n396), .A2(new_n403), .A3(new_n404), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT31), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT69), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(G472), .A2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT32), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n411), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n412), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT69), .B1(new_n412), .B2(KEYINPUT31), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT32), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n418), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n408), .A2(new_n409), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n427), .B2(new_n403), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n396), .A2(new_n404), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n402), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n384), .A2(new_n389), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n328), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT71), .A3(new_n404), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n435), .A3(new_n328), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(KEYINPUT28), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n404), .A2(new_n407), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(KEYINPUT29), .A3(new_n403), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n439), .B2(KEYINPUT72), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n431), .B(new_n440), .C1(KEYINPUT72), .C2(new_n439), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n420), .A2(new_n426), .B1(G472), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G217), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(G234), .B2(new_n191), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT25), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT22), .B(G137), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n312), .B2(G128), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n452), .B(new_n453), .C1(G119), .C2(new_n258), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G110), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G125), .B(G140), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT16), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT16), .ZN(new_n460));
  INV_X1    g274(.A(G140), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G125), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(G146), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT74), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n459), .A2(KEYINPUT74), .A3(new_n462), .A4(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n192), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT24), .B(G110), .Z(new_n470));
  XNOR2_X1  g284(.A(G119), .B(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n457), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  OAI22_X1  g287(.A1(new_n454), .A2(G110), .B1(new_n471), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n458), .A2(new_n192), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n463), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n450), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n473), .B2(new_n476), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n478), .A3(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n477), .B1(new_n482), .B2(new_n450), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n446), .B1(new_n483), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n481), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n450), .B1(new_n485), .B2(new_n479), .ZN(new_n486));
  INV_X1    g300(.A(new_n477), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n445), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n444), .A2(G902), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT76), .B1(new_n442), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n441), .A2(G472), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n417), .A2(KEYINPUT32), .A3(new_n419), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n425), .B1(new_n424), .B2(new_n418), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT76), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n492), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n469), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n398), .A2(G214), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT88), .A3(new_n194), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n194), .A2(KEYINPUT88), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(G214), .A3(new_n398), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT17), .A3(G131), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(G131), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n502), .B(new_n508), .C1(KEYINPUT17), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(KEYINPUT18), .A3(G131), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n458), .B(new_n192), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT18), .A2(G131), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n504), .A2(new_n513), .A3(new_n506), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n214), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n191), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n519), .B1(new_n510), .B2(new_n515), .ZN(new_n522));
  OAI21_X1  g336(.A(G475), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n458), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT19), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n509), .B(new_n463), .C1(G146), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n518), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n527), .A2(new_n528), .A3(new_n515), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n516), .B2(new_n518), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NOR2_X1   g345(.A1(G475), .A2(G902), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n523), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(G234), .A2(G237), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(G952), .A3(new_n275), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n537), .B(KEYINPUT92), .Z(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(G902), .A3(G953), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT21), .B(G898), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G128), .B(G143), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT13), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n258), .A2(KEYINPUT13), .A3(G143), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n237), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n544), .A2(new_n546), .B1(new_n248), .B2(new_n543), .ZN(new_n547));
  INV_X1    g361(.A(G122), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G116), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT91), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n314), .A2(G122), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n211), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n550), .A2(new_n211), .A3(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n547), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  INV_X1    g370(.A(new_n550), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n551), .B(KEYINPUT14), .ZN(new_n558));
  OAI21_X1  g372(.A(G107), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n248), .B(new_n543), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n304), .A2(new_n443), .A3(G953), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n555), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n555), .B2(new_n561), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n191), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n535), .A2(new_n542), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n381), .A2(new_n501), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n424), .B2(new_n191), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n417), .A2(new_n419), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n310), .A2(new_n492), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT93), .Z(new_n577));
  INV_X1    g391(.A(new_n187), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n579));
  INV_X1    g393(.A(new_n311), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n581), .B2(new_n378), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n566), .A2(new_n191), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n565), .B2(G478), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n563), .A2(new_n564), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT33), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n585), .B1(new_n587), .B2(G478), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n535), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n542), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n577), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT34), .B(G104), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G6));
  OAI211_X1 g407(.A(new_n568), .B(new_n523), .C1(new_n533), .C2(new_n534), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n542), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n577), .A2(new_n582), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT94), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G107), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  NAND2_X1  g413(.A1(new_n484), .A2(new_n489), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n444), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  OAI22_X1  g416(.A1(new_n485), .A2(new_n479), .B1(KEYINPUT36), .B2(new_n450), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n480), .A2(new_n481), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n606), .A2(new_n607), .A3(new_n491), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n606), .B2(new_n491), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n601), .A2(new_n602), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n609), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(new_n607), .A3(new_n491), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT96), .B1(new_n614), .B2(new_n490), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n616), .A2(new_n575), .A3(new_n569), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n381), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT37), .B(G110), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  NAND2_X1  g434(.A1(new_n581), .A2(new_n378), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n187), .A3(new_n310), .ZN(new_n622));
  INV_X1    g436(.A(G900), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n539), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n538), .A2(new_n624), .ZN(new_n625));
  OR3_X1    g439(.A1(new_n594), .A2(KEYINPUT97), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT97), .B1(new_n594), .B2(new_n625), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n498), .A2(new_n629), .A3(new_n616), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n258), .ZN(G30));
  XOR2_X1   g446(.A(new_n621), .B(KEYINPUT38), .Z(new_n633));
  NAND2_X1  g447(.A1(new_n420), .A2(new_n426), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n434), .A2(new_n402), .A3(new_n436), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n412), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n572), .B1(new_n639), .B2(new_n191), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT99), .B1(new_n634), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n644), .B(new_n640), .C1(new_n420), .C2(new_n426), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n633), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n625), .B(KEYINPUT39), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n310), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n614), .A2(new_n490), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n535), .A2(new_n568), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n654), .A2(new_n187), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n649), .A2(new_n652), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  INV_X1    g472(.A(new_n625), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n611), .A2(new_n615), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n589), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n622), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n192), .ZN(G48));
  NAND3_X1  g479(.A1(new_n621), .A2(new_n187), .A3(new_n590), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n288), .A2(new_n291), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n190), .B1(new_n667), .B2(new_n191), .ZN(new_n668));
  INV_X1    g482(.A(new_n292), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n306), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n498), .A2(new_n492), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT41), .B(G113), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND3_X1  g488(.A1(new_n621), .A2(new_n187), .A3(new_n595), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n314), .ZN(G18));
  NAND3_X1  g491(.A1(new_n498), .A2(new_n569), .A3(new_n616), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n670), .B(new_n187), .C1(new_n375), .C2(new_n379), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT100), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n582), .A2(new_n681), .A3(new_n670), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n678), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n312), .ZN(G21));
  AOI21_X1  g498(.A(new_n403), .B1(new_n437), .B2(new_n438), .ZN(new_n685));
  INV_X1    g499(.A(new_n412), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(new_n405), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n419), .B1(new_n687), .B2(new_n413), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n493), .A2(new_n573), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n542), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n670), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n187), .B(new_n655), .C1(new_n375), .C2(new_n379), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n582), .A2(KEYINPUT101), .A3(new_n655), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n548), .ZN(G24));
  NAND2_X1  g511(.A1(new_n680), .A2(new_n682), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n573), .A2(new_n688), .ZN(new_n699));
  INV_X1    g513(.A(new_n654), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n589), .A2(new_n625), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  AND3_X1   g519(.A1(new_n581), .A2(new_n378), .A3(new_n187), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n442), .A2(new_n493), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n302), .A2(new_n307), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n707), .A3(new_n709), .A4(new_n701), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n581), .A2(new_n378), .A3(new_n187), .A4(new_n709), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n498), .A2(new_n492), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  NAND4_X1  g532(.A1(new_n706), .A2(new_n707), .A3(new_n709), .A4(new_n629), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT102), .B(G134), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G36));
  AOI22_X1  g535(.A1(new_n295), .A2(new_n277), .B1(new_n297), .B2(new_n290), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT45), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n725));
  OAI221_X1 g539(.A(G469), .B1(KEYINPUT45), .B2(new_n722), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(new_n301), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n301), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n292), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n307), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n588), .ZN(new_n733));
  OR2_X1    g547(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n734));
  NAND2_X1  g548(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n535), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n733), .A2(new_n535), .ZN(new_n737));
  INV_X1    g551(.A(new_n735), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  OR3_X1    g554(.A1(new_n740), .A2(new_n575), .A3(new_n654), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n706), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n732), .A2(new_n650), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  XNOR2_X1  g560(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n731), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n730), .A2(new_n307), .A3(new_n747), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n706), .A2(new_n442), .A3(new_n493), .A4(new_n701), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n461), .ZN(G42));
  AND4_X1   g568(.A1(new_n492), .A2(new_n189), .A3(new_n307), .A4(new_n737), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n668), .A2(new_n669), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT106), .Z(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n648), .A3(new_n633), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n581), .A2(new_n378), .A3(new_n187), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n740), .A2(new_n538), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n689), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n757), .A2(new_n307), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n763), .B(new_n765), .C1(new_n751), .C2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n670), .B(new_n578), .C1(KEYINPUT112), .C2(KEYINPUT50), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n633), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n764), .A2(new_n706), .A3(new_n670), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n775), .A2(new_n573), .A3(new_n654), .A4(new_n688), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n706), .A2(new_n670), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n647), .A2(new_n777), .A3(new_n493), .A4(new_n538), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n535), .A2(new_n588), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n769), .A2(new_n774), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  INV_X1    g596(.A(new_n774), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n768), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n775), .A2(new_n714), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT114), .Z(new_n788));
  OR3_X1    g602(.A1(new_n788), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n275), .A2(G952), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n765), .B1(new_n680), .B2(new_n682), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n792), .B(new_n793), .C1(new_n778), .C2(new_n662), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n789), .A2(KEYINPUT116), .A3(new_n791), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n768), .A2(new_n783), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n782), .A3(KEYINPUT51), .A4(new_n780), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n786), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n590), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n188), .B(new_n803), .C1(new_n581), .C2(new_n378), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n381), .A2(new_n617), .B1(new_n804), .B2(new_n576), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n594), .B(KEYINPUT107), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n542), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n189), .B(new_n807), .C1(new_n375), .C2(new_n379), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n621), .A2(KEYINPUT108), .A3(new_n189), .A4(new_n807), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n576), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n805), .A2(new_n812), .A3(new_n570), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n611), .A2(new_n615), .A3(new_n659), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n535), .A2(new_n568), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n498), .A2(new_n310), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n817), .A2(new_n763), .B1(new_n713), .B2(new_n702), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n713), .A2(new_n714), .A3(new_n628), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n706), .A2(new_n703), .A3(new_n709), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n308), .A2(new_n309), .A3(new_n568), .A4(new_n535), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n706), .A2(new_n661), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n719), .A2(new_n821), .A3(new_n823), .A4(KEYINPUT109), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n813), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n671), .B1(new_n666), .B2(new_n675), .ZN(new_n827));
  INV_X1    g641(.A(new_n678), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n698), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n696), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n717), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n622), .B1(new_n663), .B2(new_n630), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n698), .B2(new_n703), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n700), .A2(new_n708), .A3(new_n625), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n642), .B2(new_n645), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n835), .B(new_n837), .C1(new_n694), .C2(new_n695), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n694), .A2(new_n695), .ZN(new_n839));
  INV_X1    g653(.A(new_n837), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT110), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n834), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n834), .C1(new_n838), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n832), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n843), .A2(new_n845), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n683), .A2(new_n696), .A3(new_n827), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT111), .B1(new_n851), .B2(new_n717), .ZN(new_n852));
  AND4_X1   g666(.A1(KEYINPUT111), .A2(new_n829), .A3(new_n830), .A4(new_n717), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n813), .A2(new_n825), .A3(KEYINPUT53), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n850), .A2(new_n855), .B1(new_n846), .B2(new_n847), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n802), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n762), .B1(new_n860), .B2(new_n861), .ZN(G75));
  NOR2_X1   g676(.A1(new_n275), .A2(G952), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n852), .A2(new_n854), .ZN(new_n865));
  INV_X1    g679(.A(new_n853), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n843), .A3(new_n845), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n846), .A2(new_n847), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n191), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n869), .B2(G210), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n356), .B(new_n351), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT55), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n864), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n867), .A2(new_n868), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(G210), .A4(G902), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n869), .B2(G210), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT118), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(G210), .A3(G902), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n876), .A4(new_n878), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n873), .B1(new_n881), .B2(new_n885), .ZN(G51));
  XNOR2_X1  g700(.A(new_n856), .B(KEYINPUT54), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n300), .B(KEYINPUT57), .Z(new_n888));
  OAI21_X1  g702(.A(new_n667), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n869), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(new_n726), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n863), .B1(new_n889), .B2(new_n891), .ZN(G54));
  INV_X1    g706(.A(new_n530), .ZN(new_n893));
  NAND2_X1  g707(.A1(KEYINPUT58), .A2(G475), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT119), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n864), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n890), .A2(new_n893), .A3(new_n895), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(G60));
  XNOR2_X1  g713(.A(new_n587), .B(KEYINPUT120), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n583), .B(KEYINPUT59), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n864), .B1(new_n887), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n859), .B2(new_n901), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(G63));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT60), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n867), .B2(new_n868), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n863), .B1(new_n909), .B2(new_n606), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n483), .B1(new_n856), .B2(new_n908), .ZN(new_n911));
  AOI211_X1 g725(.A(KEYINPUT121), .B(new_n906), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n908), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n874), .A2(new_n606), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n914), .A3(new_n864), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT61), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n912), .A2(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n540), .B2(new_n349), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n851), .A2(new_n813), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n921), .B2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n346), .B1(G898), .B2(new_n275), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G69));
  OAI21_X1  g738(.A(new_n390), .B1(new_n395), .B2(KEYINPUT30), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n526), .B(KEYINPUT122), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n651), .B1(new_n589), .B2(new_n806), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n501), .A3(new_n706), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n745), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n753), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n657), .A2(new_n834), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n932), .A2(new_n934), .A3(new_n938), .A4(new_n935), .ZN(new_n939));
  AOI211_X1 g753(.A(G953), .B(new_n928), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n928), .B1(G227), .B2(new_n275), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n707), .A2(new_n732), .A3(new_n650), .A4(new_n839), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n753), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n717), .A2(new_n719), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT125), .Z(new_n945));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n745), .A2(new_n946), .A3(new_n834), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n745), .B2(new_n834), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n943), .B(new_n945), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n941), .B1(new_n950), .B2(new_n275), .ZN(new_n951));
  OAI21_X1  g765(.A(G900), .B1(new_n928), .B2(G227), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(G953), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n940), .A2(new_n951), .A3(new_n953), .ZN(G72));
  XNOR2_X1  g768(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n572), .A2(new_n191), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n950), .B2(new_n920), .ZN(new_n958));
  INV_X1    g772(.A(new_n429), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n402), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n864), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n429), .A2(new_n403), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n937), .A2(new_n921), .A3(new_n939), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n957), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n686), .A2(KEYINPUT127), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n430), .Z(new_n966));
  AND3_X1   g780(.A1(new_n848), .A2(new_n957), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n961), .A2(new_n964), .A3(new_n967), .ZN(G57));
endmodule


