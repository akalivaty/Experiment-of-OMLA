

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  NOR2_X1 U323 ( .A1(n434), .A2(n433), .ZN(n490) );
  XNOR2_X1 U324 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n451) );
  XOR2_X1 U325 ( .A(KEYINPUT28), .B(n560), .Z(n532) );
  XOR2_X1 U326 ( .A(KEYINPUT17), .B(KEYINPUT80), .Z(n291) );
  XOR2_X1 U327 ( .A(KEYINPUT103), .B(n435), .Z(n292) );
  INV_X1 U328 ( .A(KEYINPUT45), .ZN(n459) );
  XNOR2_X1 U329 ( .A(n459), .B(KEYINPUT65), .ZN(n460) );
  XNOR2_X1 U330 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n398) );
  XNOR2_X1 U331 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U332 ( .A(n399), .B(n398), .ZN(n404) );
  INV_X1 U333 ( .A(KEYINPUT118), .ZN(n473) );
  XNOR2_X1 U334 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  INV_X1 U335 ( .A(G218GAT), .ZN(n370) );
  XNOR2_X1 U336 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U337 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U338 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U339 ( .A(n373), .B(n372), .ZN(n376) );
  XNOR2_X1 U340 ( .A(n447), .B(n446), .ZN(n450) );
  INV_X1 U341 ( .A(KEYINPUT124), .ZN(n481) );
  XNOR2_X1 U342 ( .A(n310), .B(n309), .ZN(n563) );
  XNOR2_X1 U343 ( .A(n378), .B(n377), .ZN(n523) );
  XNOR2_X1 U344 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U345 ( .A(n456), .B(G43GAT), .ZN(n457) );
  XNOR2_X1 U346 ( .A(n484), .B(n483), .ZN(G1352GAT) );
  XNOR2_X1 U347 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(G183GAT), .B(KEYINPUT81), .Z(n294) );
  XNOR2_X1 U349 ( .A(G15GAT), .B(G113GAT), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U351 ( .A(n295), .B(G99GAT), .Z(n297) );
  XOR2_X1 U352 ( .A(KEYINPUT0), .B(G127GAT), .Z(n417) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(n417), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U355 ( .A(G190GAT), .B(G134GAT), .Z(n441) );
  XNOR2_X1 U356 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n291), .B(n298), .ZN(n366) );
  XOR2_X1 U358 ( .A(n441), .B(n366), .Z(n300) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U361 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT79), .B(G120GAT), .Z(n304) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G176GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U365 ( .A(G71GAT), .B(KEYINPUT78), .Z(n306) );
  XNOR2_X1 U366 ( .A(KEYINPUT20), .B(KEYINPUT77), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U369 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n312) );
  NAND2_X1 U370 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U372 ( .A(n313), .B(KEYINPUT32), .Z(n315) );
  XOR2_X1 U373 ( .A(G120GAT), .B(G57GAT), .Z(n416) );
  XOR2_X1 U374 ( .A(G176GAT), .B(G64GAT), .Z(n369) );
  XNOR2_X1 U375 ( .A(n416), .B(n369), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n317) );
  XNOR2_X1 U377 ( .A(G71GAT), .B(KEYINPUT69), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n316), .B(KEYINPUT13), .ZN(n344) );
  XOR2_X1 U379 ( .A(n317), .B(n344), .Z(n323) );
  XOR2_X1 U380 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n392) );
  XOR2_X1 U383 ( .A(KEYINPUT70), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n439) );
  XNOR2_X1 U386 ( .A(n392), .B(n439), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n580) );
  XOR2_X1 U388 ( .A(G29GAT), .B(KEYINPUT8), .Z(n325) );
  XNOR2_X1 U389 ( .A(G43GAT), .B(G36GAT), .ZN(n324) );
  XNOR2_X1 U390 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U391 ( .A(G50GAT), .B(KEYINPUT7), .Z(n326) );
  XOR2_X1 U392 ( .A(n327), .B(n326), .Z(n448) );
  XOR2_X1 U393 ( .A(G113GAT), .B(G1GAT), .Z(n423) );
  XOR2_X1 U394 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n329) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U397 ( .A(n423), .B(n330), .Z(n331) );
  XOR2_X1 U398 ( .A(n448), .B(n331), .Z(n335) );
  XOR2_X1 U399 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n333) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(G141GAT), .ZN(n332) );
  XNOR2_X1 U401 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U402 ( .A(n335), .B(n334), .Z(n337) );
  XOR2_X1 U403 ( .A(G169GAT), .B(G8GAT), .Z(n374) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G15GAT), .Z(n341) );
  XNOR2_X1 U405 ( .A(n374), .B(n341), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n337), .B(n336), .ZN(n546) );
  XNOR2_X1 U407 ( .A(KEYINPUT68), .B(n546), .ZN(n564) );
  NOR2_X1 U408 ( .A1(n580), .A2(n564), .ZN(n491) );
  XOR2_X1 U409 ( .A(G78GAT), .B(G211GAT), .Z(n339) );
  XNOR2_X1 U410 ( .A(G127GAT), .B(G155GAT), .ZN(n338) );
  XNOR2_X1 U411 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U412 ( .A(n340), .B(G57GAT), .Z(n343) );
  XNOR2_X1 U413 ( .A(n341), .B(G1GAT), .ZN(n342) );
  XNOR2_X1 U414 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U415 ( .A(G183GAT), .B(KEYINPUT73), .Z(n368) );
  XOR2_X1 U416 ( .A(n368), .B(n344), .Z(n346) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U419 ( .A(n348), .B(n347), .Z(n356) );
  XOR2_X1 U420 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n350) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(G64GAT), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT74), .Z(n352) );
  XNOR2_X1 U424 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U427 ( .A(n356), .B(n355), .Z(n553) );
  INV_X1 U428 ( .A(n553), .ZN(n584) );
  XOR2_X1 U429 ( .A(KEYINPUT92), .B(G92GAT), .Z(n358) );
  XNOR2_X1 U430 ( .A(G190GAT), .B(G204GAT), .ZN(n357) );
  XOR2_X1 U431 ( .A(n358), .B(n357), .Z(n378) );
  XNOR2_X1 U432 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n359), .B(G211GAT), .ZN(n393) );
  INV_X1 U434 ( .A(n393), .ZN(n361) );
  INV_X1 U435 ( .A(KEYINPUT93), .ZN(n360) );
  NAND2_X1 U436 ( .A1(n361), .A2(n360), .ZN(n363) );
  NAND2_X1 U437 ( .A1(n393), .A2(KEYINPUT93), .ZN(n362) );
  NAND2_X1 U438 ( .A1(n363), .A2(n362), .ZN(n365) );
  AND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U440 ( .A(n365), .B(n364), .ZN(n367) );
  XNOR2_X1 U441 ( .A(n367), .B(n366), .ZN(n373) );
  XOR2_X1 U442 ( .A(n369), .B(n368), .Z(n371) );
  XNOR2_X1 U443 ( .A(G36GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  NOR2_X1 U445 ( .A1(n563), .A2(n523), .ZN(n397) );
  XNOR2_X1 U446 ( .A(G155GAT), .B(KEYINPUT84), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n379), .B(KEYINPUT3), .ZN(n380) );
  XOR2_X1 U448 ( .A(n380), .B(KEYINPUT2), .Z(n382) );
  XNOR2_X1 U449 ( .A(G141GAT), .B(G162GAT), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n422) );
  XOR2_X1 U451 ( .A(G218GAT), .B(KEYINPUT71), .Z(n440) );
  XOR2_X1 U452 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n384) );
  XNOR2_X1 U453 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U455 ( .A(n440), .B(n385), .Z(n387) );
  NAND2_X1 U456 ( .A1(G228GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U457 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U458 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n389) );
  XNOR2_X1 U459 ( .A(G22GAT), .B(KEYINPUT85), .ZN(n388) );
  XNOR2_X1 U460 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U461 ( .A(n391), .B(n390), .Z(n395) );
  XNOR2_X1 U462 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n422), .B(n396), .ZN(n560) );
  NOR2_X1 U465 ( .A1(n397), .A2(n560), .ZN(n399) );
  NAND2_X1 U466 ( .A1(n560), .A2(n563), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n400), .B(KEYINPUT26), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n401), .B(KEYINPUT96), .ZN(n545) );
  XOR2_X1 U469 ( .A(KEYINPUT27), .B(KEYINPUT94), .Z(n402) );
  XOR2_X1 U470 ( .A(n523), .B(n402), .Z(n429) );
  NOR2_X1 U471 ( .A1(n545), .A2(n429), .ZN(n403) );
  NOR2_X1 U472 ( .A1(n404), .A2(n403), .ZN(n426) );
  XOR2_X1 U473 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n406) );
  XNOR2_X1 U474 ( .A(G134GAT), .B(G148GAT), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U476 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT1), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U479 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U480 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n412) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U482 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U483 ( .A(KEYINPUT5), .B(n413), .ZN(n414) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U485 ( .A(G85GAT), .B(n416), .Z(n419) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U488 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n428) );
  NOR2_X1 U491 ( .A1(n426), .A2(n428), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n427), .B(KEYINPUT98), .ZN(n434) );
  INV_X1 U493 ( .A(n532), .ZN(n432) );
  XNOR2_X1 U494 ( .A(KEYINPUT91), .B(n428), .ZN(n521) );
  NOR2_X1 U495 ( .A1(n429), .A2(n521), .ZN(n430) );
  XOR2_X1 U496 ( .A(KEYINPUT95), .B(n430), .Z(n530) );
  NAND2_X1 U497 ( .A1(n530), .A2(n563), .ZN(n431) );
  NOR2_X1 U498 ( .A1(n432), .A2(n431), .ZN(n433) );
  NOR2_X1 U499 ( .A1(n584), .A2(n490), .ZN(n435) );
  XOR2_X1 U500 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n437) );
  XNOR2_X1 U501 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n436) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U503 ( .A(n439), .B(n438), .Z(n447) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U505 ( .A(G106GAT), .B(KEYINPUT72), .Z(n443) );
  NAND2_X1 U506 ( .A1(G232GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n448), .B(G162GAT), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n575) );
  XNOR2_X1 U510 ( .A(KEYINPUT36), .B(n575), .ZN(n586) );
  NAND2_X1 U511 ( .A1(n292), .A2(n586), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n519) );
  NAND2_X1 U513 ( .A1(n491), .A2(n519), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT38), .B(KEYINPUT105), .Z(n453) );
  XNOR2_X1 U515 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U516 ( .A(KEYINPUT106), .B(n455), .ZN(n506) );
  NOR2_X1 U517 ( .A1(n563), .A2(n506), .ZN(n458) );
  INV_X1 U518 ( .A(KEYINPUT40), .ZN(n456) );
  INV_X1 U519 ( .A(n523), .ZN(n472) );
  NAND2_X1 U520 ( .A1(n584), .A2(n586), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n580), .A2(n462), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n463), .A2(n564), .ZN(n470) );
  XOR2_X1 U523 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n468) );
  XNOR2_X1 U524 ( .A(n580), .B(KEYINPUT41), .ZN(n550) );
  NOR2_X1 U525 ( .A1(n546), .A2(n550), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n464), .B(KEYINPUT46), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n584), .A2(n465), .ZN(n466) );
  INV_X1 U528 ( .A(n575), .ZN(n557) );
  NAND2_X1 U529 ( .A1(n466), .A2(n557), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT48), .ZN(n531) );
  NAND2_X1 U533 ( .A1(n472), .A2(n531), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n476), .A2(n521), .ZN(n559) );
  NOR2_X1 U535 ( .A1(n545), .A2(n559), .ZN(n477) );
  XOR2_X1 U536 ( .A(n477), .B(KEYINPUT123), .Z(n587) );
  INV_X1 U537 ( .A(n587), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n546), .A2(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n484) );
  XNOR2_X1 U541 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n482) );
  NOR2_X1 U542 ( .A1(n506), .A2(n523), .ZN(n487) );
  INV_X1 U543 ( .A(G36GAT), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(KEYINPUT108), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  NOR2_X1 U546 ( .A1(n575), .A2(n553), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n488), .Z(n489) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n508) );
  NAND2_X1 U549 ( .A1(n491), .A2(n508), .ZN(n500) );
  NOR2_X1 U550 ( .A1(n521), .A2(n500), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(n492), .Z(n493) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n523), .A2(n500), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(n496), .ZN(G1325GAT) );
  NOR2_X1 U557 ( .A1(n563), .A2(n500), .ZN(n498) );
  XNOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U560 ( .A(G15GAT), .B(n499), .Z(G1326GAT) );
  NOR2_X1 U561 ( .A1(n532), .A2(n500), .ZN(n501) );
  XOR2_X1 U562 ( .A(G22GAT), .B(n501), .Z(G1327GAT) );
  NOR2_X1 U563 ( .A1(n506), .A2(n521), .ZN(n505) );
  XOR2_X1 U564 ( .A(KEYINPUT102), .B(KEYINPUT107), .Z(n503) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n532), .A2(n506), .ZN(n507) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT109), .B(n550), .ZN(n568) );
  AND2_X1 U571 ( .A1(n546), .A2(n568), .ZN(n520) );
  NAND2_X1 U572 ( .A1(n520), .A2(n508), .ZN(n516) );
  NOR2_X1 U573 ( .A1(n521), .A2(n516), .ZN(n509) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n516), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n563), .A2(n516), .ZN(n514) );
  XOR2_X1 U581 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n532), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U587 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n527), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U592 ( .A1(n563), .A2(n527), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n532), .A2(n527), .ZN(n528) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n544) );
  NOR2_X1 U598 ( .A1(n563), .A2(n544), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n535) );
  NOR2_X1 U600 ( .A1(n564), .A2(n535), .ZN(n534) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  INV_X1 U603 ( .A(n535), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n541), .A2(n568), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U607 ( .A1(n541), .A2(n584), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U611 ( .A1(n541), .A2(n575), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  OR2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n546), .A2(n556), .ZN(n547) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n550), .A2(n556), .ZN(n551) );
  XOR2_X1 U620 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NOR2_X1 U621 ( .A1(n553), .A2(n556), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT119), .Z(n567) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT55), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n576) );
  INV_X1 U630 ( .A(n564), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n572) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT120), .Z(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n576), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  XOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT121), .Z(n574) );
  NAND2_X1 U639 ( .A1(n576), .A2(n584), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G190GAT), .B(n579), .Z(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U646 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

