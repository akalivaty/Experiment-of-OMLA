

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U323 ( .A(G92GAT), .B(G85GAT), .Z(n367) );
  XNOR2_X1 U324 ( .A(n383), .B(n382), .ZN(n389) );
  XNOR2_X1 U325 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U326 ( .A(n375), .B(n291), .ZN(n376) );
  XOR2_X1 U327 ( .A(n374), .B(n373), .Z(n291) );
  XNOR2_X1 U328 ( .A(n381), .B(KEYINPUT47), .ZN(n382) );
  XOR2_X1 U329 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  INV_X1 U330 ( .A(KEYINPUT48), .ZN(n390) );
  XNOR2_X1 U331 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U332 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U333 ( .A(n344), .B(n343), .ZN(n385) );
  INV_X1 U334 ( .A(G183GAT), .ZN(n458) );
  XNOR2_X1 U335 ( .A(n455), .B(G190GAT), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n435) );
  XOR2_X1 U338 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n293) );
  XNOR2_X1 U339 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n311) );
  XOR2_X1 U341 ( .A(G162GAT), .B(G57GAT), .Z(n295) );
  XNOR2_X1 U342 ( .A(G134GAT), .B(G127GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U344 ( .A(G148GAT), .B(G120GAT), .Z(n297) );
  XNOR2_X1 U345 ( .A(G1GAT), .B(G141GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U347 ( .A(n299), .B(n298), .Z(n305) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n300), .B(KEYINPUT83), .ZN(n447) );
  XOR2_X1 U350 ( .A(G85GAT), .B(n447), .Z(n302) );
  NAND2_X1 U351 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U355 ( .A(n306), .B(KEYINPUT93), .Z(n309) );
  XNOR2_X1 U356 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n307), .B(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U358 ( .A(n420), .B(KEYINPUT94), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U360 ( .A(n311), .B(n310), .Z(n505) );
  INV_X1 U361 ( .A(n505), .ZN(n520) );
  XOR2_X1 U362 ( .A(G8GAT), .B(KEYINPUT79), .Z(n400) );
  XOR2_X1 U363 ( .A(n400), .B(G64GAT), .Z(n313) );
  XOR2_X1 U364 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XNOR2_X1 U365 ( .A(n439), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n314), .B(KEYINPUT14), .Z(n320) );
  XNOR2_X1 U368 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n315), .B(KEYINPUT73), .ZN(n338) );
  XOR2_X1 U370 ( .A(G78GAT), .B(n338), .Z(n317) );
  NAND2_X1 U371 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U373 ( .A(G183GAT), .B(n318), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U375 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n322) );
  XNOR2_X1 U376 ( .A(G22GAT), .B(KEYINPUT12), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U378 ( .A(KEYINPUT81), .B(G155GAT), .Z(n324) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U381 ( .A(n326), .B(n325), .Z(n327) );
  XOR2_X1 U382 ( .A(n328), .B(n327), .Z(n579) );
  INV_X1 U383 ( .A(n579), .ZN(n555) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G71GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n329), .B(G120GAT), .ZN(n449) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(n449), .ZN(n331) );
  XOR2_X1 U387 ( .A(KEYINPUT32), .B(n367), .Z(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U389 ( .A(G64GAT), .B(KEYINPUT75), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n332), .B(G204GAT), .ZN(n399) );
  XOR2_X1 U391 ( .A(n399), .B(KEYINPUT76), .Z(n334) );
  NAND2_X1 U392 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U394 ( .A(n336), .B(n335), .Z(n344) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(G78GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n337), .B(G148GAT), .ZN(n421) );
  XNOR2_X1 U397 ( .A(n338), .B(n421), .ZN(n342) );
  XOR2_X1 U398 ( .A(KEYINPUT77), .B(KEYINPUT74), .Z(n340) );
  XNOR2_X1 U399 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n339) );
  XOR2_X1 U400 ( .A(n340), .B(n339), .Z(n341) );
  XOR2_X1 U401 ( .A(KEYINPUT41), .B(KEYINPUT65), .Z(n345) );
  XOR2_X1 U402 ( .A(n385), .B(n345), .Z(n561) );
  XOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT72), .Z(n347) );
  XNOR2_X1 U404 ( .A(G1GAT), .B(G113GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n363) );
  XOR2_X1 U406 ( .A(G197GAT), .B(G8GAT), .Z(n349) );
  XNOR2_X1 U407 ( .A(G50GAT), .B(G43GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U409 ( .A(n350), .B(G15GAT), .Z(n352) );
  XOR2_X1 U410 ( .A(G22GAT), .B(G141GAT), .Z(n429) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(n429), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U413 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n354) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U416 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U417 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n358) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G29GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U420 ( .A(KEYINPUT8), .B(n359), .Z(n379) );
  XNOR2_X1 U421 ( .A(n379), .B(KEYINPUT29), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n569) );
  OR2_X1 U424 ( .A1(n561), .A2(n569), .ZN(n365) );
  XNOR2_X1 U425 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  NOR2_X1 U427 ( .A1(n555), .A2(n366), .ZN(n380) );
  XOR2_X1 U428 ( .A(n367), .B(n428), .Z(n369) );
  NAND2_X1 U429 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n377) );
  XOR2_X1 U431 ( .A(G43GAT), .B(G134GAT), .Z(n440) );
  XOR2_X1 U432 ( .A(KEYINPUT11), .B(KEYINPUT67), .Z(n371) );
  XNOR2_X1 U433 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n440), .B(n372), .ZN(n375) );
  XOR2_X1 U436 ( .A(KEYINPUT10), .B(G106GAT), .Z(n374) );
  XNOR2_X1 U437 ( .A(G190GAT), .B(G99GAT), .ZN(n373) );
  XOR2_X1 U438 ( .A(n379), .B(n378), .Z(n557) );
  INV_X1 U439 ( .A(n557), .ZN(n473) );
  NAND2_X1 U440 ( .A1(n380), .A2(n473), .ZN(n383) );
  XOR2_X1 U441 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n381) );
  XOR2_X1 U442 ( .A(KEYINPUT36), .B(n557), .Z(n582) );
  NOR2_X1 U443 ( .A1(n582), .A2(n579), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n384), .B(KEYINPUT45), .ZN(n386) );
  BUF_X1 U445 ( .A(n385), .Z(n575) );
  NAND2_X1 U446 ( .A1(n386), .A2(n575), .ZN(n387) );
  INV_X1 U447 ( .A(n569), .ZN(n549) );
  NOR2_X1 U448 ( .A1(n387), .A2(n549), .ZN(n388) );
  NOR2_X1 U449 ( .A1(n389), .A2(n388), .ZN(n393) );
  XOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT112), .Z(n391) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n548) );
  INV_X1 U452 ( .A(n548), .ZN(n530) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n395) );
  XNOR2_X1 U454 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U456 ( .A(n396), .B(G183GAT), .Z(n398) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(G176GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n450) );
  XOR2_X1 U459 ( .A(n400), .B(n399), .Z(n402) );
  XNOR2_X1 U460 ( .A(G36GAT), .B(G92GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U462 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n404) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U465 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U466 ( .A(KEYINPUT91), .B(G218GAT), .Z(n408) );
  XNOR2_X1 U467 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U469 ( .A(G197GAT), .B(n409), .ZN(n432) );
  XOR2_X1 U470 ( .A(n432), .B(KEYINPUT97), .Z(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n450), .B(n412), .ZN(n508) );
  INV_X1 U473 ( .A(n508), .ZN(n522) );
  NAND2_X1 U474 ( .A1(n530), .A2(n522), .ZN(n414) );
  XOR2_X1 U475 ( .A(KEYINPUT54), .B(KEYINPUT117), .Z(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U477 ( .A1(n520), .A2(n415), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n416), .B(KEYINPUT66), .ZN(n568) );
  XOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n418) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U482 ( .A(n419), .B(KEYINPUT92), .Z(n423) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n425) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT89), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U488 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n464) );
  NAND2_X1 U492 ( .A1(n568), .A2(n464), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U494 ( .A(KEYINPUT55), .B(n436), .ZN(n453) );
  XOR2_X1 U495 ( .A(KEYINPUT84), .B(KEYINPUT87), .Z(n438) );
  XNOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT86), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n442) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U504 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U506 ( .A(n452), .B(n451), .Z(n511) );
  INV_X1 U507 ( .A(n511), .ZN(n531) );
  NAND2_X1 U508 ( .A1(n453), .A2(n531), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n454), .B(KEYINPUT120), .ZN(n562) );
  NOR2_X1 U510 ( .A1(n562), .A2(n473), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n455) );
  NOR2_X1 U512 ( .A1(n579), .A2(n562), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT122), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n460), .B(n459), .ZN(G1350GAT) );
  XOR2_X1 U515 ( .A(n508), .B(KEYINPUT27), .Z(n466) );
  AND2_X1 U516 ( .A1(n520), .A2(n466), .ZN(n546) );
  XOR2_X1 U517 ( .A(n464), .B(KEYINPUT28), .Z(n526) );
  INV_X1 U518 ( .A(n526), .ZN(n514) );
  NAND2_X1 U519 ( .A1(n546), .A2(n514), .ZN(n533) );
  XOR2_X1 U520 ( .A(KEYINPUT88), .B(n511), .Z(n461) );
  NOR2_X1 U521 ( .A1(n533), .A2(n461), .ZN(n472) );
  NAND2_X1 U522 ( .A1(n531), .A2(n522), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n464), .A2(n462), .ZN(n463) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n463), .Z(n468) );
  NOR2_X1 U525 ( .A1(n464), .A2(n531), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT26), .ZN(n567) );
  NAND2_X1 U527 ( .A1(n567), .A2(n466), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT98), .B(n469), .Z(n470) );
  NOR2_X1 U530 ( .A1(n520), .A2(n470), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n487) );
  NAND2_X1 U532 ( .A1(n555), .A2(n473), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT82), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT16), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n487), .A2(n476), .ZN(n504) );
  NAND2_X1 U536 ( .A1(n575), .A2(n549), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT78), .B(n477), .Z(n491) );
  NAND2_X1 U538 ( .A1(n504), .A2(n491), .ZN(n484) );
  NOR2_X1 U539 ( .A1(n505), .A2(n484), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n508), .A2(n484), .ZN(n481) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n511), .A2(n484), .ZN(n483) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n514), .A2(n484), .ZN(n485) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(n485), .Z(n486) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(KEYINPUT37), .Z(n490) );
  NOR2_X1 U552 ( .A1(n582), .A2(n487), .ZN(n488) );
  NAND2_X1 U553 ( .A1(n579), .A2(n488), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n517) );
  NAND2_X1 U555 ( .A1(n491), .A2(n517), .ZN(n492) );
  XOR2_X1 U556 ( .A(KEYINPUT38), .B(n492), .Z(n501) );
  NAND2_X1 U557 ( .A1(n520), .A2(n501), .ZN(n494) );
  XOR2_X1 U558 ( .A(KEYINPUT39), .B(KEYINPUT102), .Z(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(n495), .ZN(G1328GAT) );
  XOR2_X1 U561 ( .A(G36GAT), .B(KEYINPUT103), .Z(n497) );
  NAND2_X1 U562 ( .A1(n522), .A2(n501), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n499) );
  NAND2_X1 U565 ( .A1(n531), .A2(n501), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U567 ( .A(G43GAT), .B(n500), .Z(G1330GAT) );
  XOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U569 ( .A1(n526), .A2(n501), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  NOR2_X1 U571 ( .A1(n549), .A2(n561), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n518), .A2(n504), .ZN(n513) );
  NOR2_X1 U573 ( .A1(n505), .A2(n513), .ZN(n506) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n506), .Z(n507) );
  XNOR2_X1 U575 ( .A(KEYINPUT42), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U576 ( .A1(n508), .A2(n513), .ZN(n509) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(n509), .Z(n510) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U579 ( .A1(n511), .A2(n513), .ZN(n512) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(KEYINPUT107), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n527), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(KEYINPUT108), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n531), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n543), .A2(n549), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n536) );
  INV_X1 U601 ( .A(n561), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n543), .A2(n551), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n539) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n555), .A2(n543), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n540), .B(KEYINPUT114), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U612 ( .A1(n543), .A2(n557), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n546), .A2(n567), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n549), .A2(n558), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U619 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n558), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n562), .A2(n569), .ZN(n560) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n560), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n581) );
  NOR2_X1 U634 ( .A1(n569), .A2(n581), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

