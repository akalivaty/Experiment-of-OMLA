//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n541, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  AND3_X1   g035(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n464), .A2(G136), .ZN(new_n473));
  AND2_X1   g048(.A1(G112), .A2(G2105), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n474), .B1(G100), .B2(new_n470), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n458), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n461), .A2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(new_n479), .B2(G124), .ZN(G162));
  AND3_X1   g055(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .ZN(new_n481));
  AND2_X1   g056(.A1(G102), .A2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n470), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(G114), .A2(G2104), .ZN(new_n484));
  INV_X1    g059(.A(G126), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n463), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n468), .A2(G138), .A3(new_n470), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n486), .A2(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G651), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(new_n496), .B1(new_n493), .B2(G651), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G88), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G50), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n505), .A2(new_n495), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(G303));
  INV_X1    g082(.A(G303), .ZN(G166));
  NAND3_X1  g083(.A1(new_n497), .A2(G89), .A3(new_n498), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT69), .B(G51), .Z(new_n510));
  NAND3_X1  g085(.A1(new_n497), .A2(G543), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(G63), .A2(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT7), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n515), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n498), .A2(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n509), .A2(new_n511), .A3(new_n517), .ZN(G168));
  NAND3_X1  g093(.A1(new_n497), .A2(G52), .A3(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n497), .A2(G90), .A3(new_n498), .ZN(new_n520));
  INV_X1    g095(.A(G64), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(G77), .A2(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(G171));
  INV_X1    g102(.A(G56), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n522), .B2(new_n523), .ZN(new_n529));
  AND2_X1   g104(.A1(G68), .A2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(G651), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n494), .A2(new_n496), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n493), .A2(G651), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n532), .A2(G43), .A3(G543), .A4(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(G81), .A3(new_n533), .A4(new_n498), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT70), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G188));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n532), .A2(G53), .A3(G543), .A4(new_n533), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT9), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n497), .A2(new_n548), .A3(G53), .A4(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AND4_X1   g125(.A1(G91), .A2(new_n532), .A3(new_n533), .A4(new_n498), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(KEYINPUT5), .A2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(KEYINPUT5), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(G65), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(KEYINPUT71), .A3(new_n556), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(G651), .A3(new_n560), .ZN(new_n561));
  AND4_X1   g136(.A1(new_n545), .A2(new_n550), .A3(new_n552), .A4(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n556), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n498), .B2(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n495), .B1(new_n564), .B2(KEYINPUT71), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n551), .B1(new_n565), .B2(new_n559), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n545), .B1(new_n566), .B2(new_n550), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  NAND3_X1  g143(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(G301));
  NAND3_X1  g144(.A1(new_n509), .A2(new_n511), .A3(new_n517), .ZN(G286));
  NAND2_X1  g145(.A1(new_n500), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n503), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n500), .A2(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n503), .A2(G48), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n498), .A2(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT73), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n503), .A2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n500), .A2(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n495), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n553), .A2(new_n554), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n502), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n500), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n499), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n596), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n589), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n589), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  XOR2_X1   g182(.A(G299), .B(KEYINPUT76), .Z(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  MUX2_X1   g188(.A(new_n536), .B(new_n613), .S(G868), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n479), .A2(G123), .ZN(new_n616));
  MUX2_X1   g191(.A(G99), .B(G111), .S(G2105), .Z(new_n617));
  AOI22_X1  g192(.A1(new_n464), .A2(G135), .B1(G2104), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G2096), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(KEYINPUT78), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(KEYINPUT78), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n624), .A2(KEYINPUT13), .ZN(new_n629));
  OR3_X1    g204(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n627), .B2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n621), .A2(new_n630), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT79), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n641), .B2(new_n643), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n638), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT80), .Z(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT17), .Z(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT81), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n654), .ZN(new_n657));
  INV_X1    g232(.A(new_n650), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n653), .C1(new_n658), .C2(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n652), .A3(new_n654), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n656), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n620), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT20), .Z(new_n673));
  AOI211_X1 g248(.A(new_n671), .B(new_n673), .C1(new_n666), .C2(new_n670), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  AND2_X1   g256(.A1(KEYINPUT24), .A2(G34), .ZN(new_n682));
  NOR2_X1   g257(.A1(KEYINPUT24), .A2(G34), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G160), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n681), .ZN(new_n686));
  INV_X1    g261(.A(G2084), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT92), .Z(new_n689));
  AND2_X1   g264(.A1(new_n479), .A2(G129), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n464), .A2(G141), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n459), .A2(G105), .ZN(new_n692));
  NAND3_X1  g267(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT26), .Z(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(new_n681), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n681), .B2(G32), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT27), .B(G1996), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n681), .A2(G33), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n468), .A2(G127), .ZN(new_n702));
  INV_X1    g277(.A(G115), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n458), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n470), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n705), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT91), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n464), .A2(G139), .ZN(new_n709));
  INV_X1    g284(.A(new_n459), .ZN(new_n710));
  INV_X1    g285(.A(G103), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT25), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR3_X1    g287(.A1(new_n710), .A2(KEYINPUT25), .A3(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT89), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n701), .B1(new_n716), .B2(new_n681), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G2072), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G2072), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n700), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n686), .A2(new_n687), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NOR2_X1   g298(.A1(G171), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G5), .B2(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(G1961), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n722), .B(new_n727), .C1(new_n698), .C2(new_n699), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT95), .Z(new_n729));
  AND2_X1   g304(.A1(KEYINPUT30), .A2(G28), .ZN(new_n730));
  NOR2_X1   g305(.A1(KEYINPUT30), .A2(G28), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n681), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT31), .B(G11), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n732), .B(new_n733), .C1(new_n619), .C2(new_n681), .ZN(new_n734));
  NAND2_X1  g309(.A1(G164), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G27), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n736), .A2(new_n737), .B1(new_n726), .B2(new_n725), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n734), .B(new_n738), .C1(new_n737), .C2(new_n736), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT94), .B1(G16), .B2(G21), .ZN(new_n740));
  NAND2_X1  g315(.A1(G168), .A2(G16), .ZN(new_n741));
  MUX2_X1   g316(.A(KEYINPUT94), .B(new_n740), .S(new_n741), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1966), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G299), .A2(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n723), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2090), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n729), .A2(new_n744), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n721), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G22), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G166), .B2(G16), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1971), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n723), .A2(G23), .ZN(new_n759));
  INV_X1    g334(.A(G288), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n723), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT33), .B(G1976), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G6), .A2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G305), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT32), .B(G1981), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  OR3_X1    g344(.A1(new_n764), .A2(KEYINPUT34), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G25), .A2(G29), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT82), .ZN(new_n772));
  INV_X1    g347(.A(G131), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n465), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n464), .A2(KEYINPUT82), .A3(G131), .ZN(new_n775));
  MUX2_X1   g350(.A(G95), .B(G107), .S(G2105), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n774), .A2(new_n775), .B1(G2104), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n479), .A2(G119), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n771), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT35), .B(G1991), .Z(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n781), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  OR2_X1    g360(.A1(G16), .A2(G24), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G290), .B2(new_n723), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT34), .B1(new_n764), .B2(new_n769), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n787), .A2(new_n785), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n770), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(KEYINPUT36), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(KEYINPUT36), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT84), .ZN(new_n798));
  INV_X1    g373(.A(new_n604), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n723), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G19), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n537), .B2(G16), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT85), .B(G1341), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n681), .A2(G26), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT28), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n464), .A2(G140), .ZN(new_n808));
  NOR2_X1   g383(.A1(G104), .A2(G2105), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT86), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n479), .B2(G128), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n681), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT87), .B(G2067), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n801), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT88), .Z(new_n818));
  NAND4_X1  g393(.A1(new_n755), .A2(new_n795), .A3(new_n796), .A4(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NAND2_X1  g395(.A1(new_n604), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n536), .A2(KEYINPUT97), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n531), .A2(new_n534), .A3(new_n535), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n497), .A2(G55), .A3(G543), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n497), .A2(G93), .A3(new_n498), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n522), .B2(new_n523), .ZN(new_n830));
  AND2_X1   g405(.A1(G80), .A2(G543), .ZN(new_n831));
  OAI21_X1  g406(.A(G651), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n824), .A2(new_n826), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n826), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n823), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  OR2_X1    g418(.A1(new_n840), .A2(new_n843), .ZN(G145));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n846), .B(new_n847), .C1(G118), .C2(new_n470), .ZN(new_n848));
  INV_X1    g423(.A(G142), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n465), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n479), .B2(G130), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n779), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n624), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT101), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n852), .B(new_n853), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n813), .B(new_n490), .ZN(new_n860));
  INV_X1    g435(.A(new_n696), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n708), .A2(new_n715), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n716), .A2(KEYINPUT99), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n865), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n868), .A2(new_n862), .A3(new_n863), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n859), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n858), .A3(new_n856), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G162), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n619), .ZN(new_n876));
  AOI21_X1  g451(.A(G37), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n872), .B2(new_n857), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n881), .B2(new_n873), .ZN(new_n882));
  INV_X1    g457(.A(new_n873), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n883), .A2(new_n880), .A3(KEYINPUT102), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n877), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g461(.A1(new_n833), .A2(G868), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n613), .B(new_n836), .Z(new_n888));
  AND2_X1   g463(.A1(new_n547), .A2(new_n549), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n560), .A2(G651), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT71), .B1(new_n555), .B2(new_n556), .ZN(new_n891));
  INV_X1    g466(.A(G91), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(new_n499), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT72), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n566), .A2(new_n545), .A3(new_n550), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n601), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n601), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT41), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n597), .A2(new_n600), .ZN(new_n900));
  INV_X1    g475(.A(new_n596), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n562), .B2(new_n567), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  OAI211_X1 g481(.A(KEYINPUT103), .B(new_n902), .C1(new_n562), .C2(new_n567), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n896), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n888), .A2(new_n899), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n897), .A2(new_n898), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n888), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  XNOR2_X1  g491(.A(G288), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(G303), .B(G305), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT106), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n915), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n887), .B1(new_n923), .B2(G868), .ZN(G295));
  AOI21_X1  g499(.A(new_n887), .B1(new_n923), .B2(G868), .ZN(G331));
  NAND2_X1  g500(.A1(G171), .A2(G168), .ZN(new_n926));
  NAND2_X1  g501(.A1(G301), .A2(G286), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n836), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n834), .A2(new_n835), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n834), .A2(new_n835), .A3(new_n927), .A4(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n908), .A2(new_n935), .A3(new_n899), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT108), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n908), .A2(new_n935), .A3(new_n938), .A4(new_n899), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n919), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n918), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n929), .A2(new_n934), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n913), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n940), .B2(new_n944), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n896), .B1(new_n898), .B2(KEYINPUT103), .ZN(new_n950));
  INV_X1    g525(.A(new_n907), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT41), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(KEYINPUT41), .A3(new_n943), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n934), .B1(new_n931), .B2(new_n932), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n836), .A2(new_n932), .A3(new_n928), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n952), .B2(new_n943), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n953), .B1(new_n957), .B2(new_n913), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n958), .B2(new_n920), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n945), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n949), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n959), .A2(new_n945), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n959), .A2(KEYINPUT110), .A3(new_n945), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n960), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n940), .A2(new_n944), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n920), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(new_n960), .A3(new_n946), .A4(new_n945), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT44), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n972), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n947), .A2(new_n948), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n966), .B1(new_n979), .B2(new_n960), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n959), .A2(KEYINPUT110), .A3(new_n945), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT110), .B1(new_n959), .B2(new_n945), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT43), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT111), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n967), .B1(new_n978), .B2(new_n984), .ZN(G397));
  AOI21_X1  g560(.A(G1384), .B1(new_n483), .B2(new_n489), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n987));
  INV_X1    g562(.A(G40), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n467), .A2(new_n988), .A3(new_n471), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n990), .A2(new_n991), .A3(new_n696), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT112), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(G1996), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n813), .B(G2067), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n995), .A2(new_n861), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n990), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n780), .A2(new_n782), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n779), .A2(new_n783), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G290), .B(G1986), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n986), .A2(new_n989), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G305), .A2(G1981), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(KEYINPUT116), .A3(new_n1014), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1012), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1019), .A2(G1976), .A3(G288), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1009), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1007), .B(KEYINPUT117), .Z(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n490), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G160), .A2(G40), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n986), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1025), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1034), .A2(new_n987), .A3(new_n1029), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1033), .A2(G2090), .B1(new_n1035), .B2(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G303), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1036), .B(G8), .C1(new_n1040), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n760), .A2(G1976), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1008), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n760), .B2(G1976), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(new_n1019), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1022), .A2(new_n1023), .B1(new_n1044), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT63), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1035), .A2(G1971), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1031), .A2(new_n1026), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G2090), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1043), .A2(new_n1040), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1051), .A2(new_n1060), .A3(new_n1044), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1028), .A2(new_n1032), .A3(new_n1031), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n687), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n987), .B2(new_n1029), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1034), .A2(KEYINPUT119), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT118), .B(new_n989), .C1(new_n986), .C2(KEYINPUT45), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1966), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1062), .B1(new_n1064), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G168), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1054), .B1(new_n1061), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1036), .A2(G8), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1054), .B1(new_n1079), .B2(new_n1059), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1080), .A3(new_n1044), .A4(new_n1051), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1053), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1035), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT120), .B(G1956), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1056), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n566), .A2(KEYINPUT57), .A3(new_n550), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(KEYINPUT122), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n550), .B1(new_n893), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n566), .A2(KEYINPUT121), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1088), .A2(KEYINPUT122), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1033), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n986), .A2(new_n989), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G2067), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1099), .A2(new_n1108), .A3(new_n604), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1035), .A2(new_n1083), .B1(new_n1056), .B2(new_n1085), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1096), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT61), .B1(new_n1110), .B2(new_n1096), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n987), .A2(new_n1029), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n991), .A3(new_n1069), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND3_X1  g691(.A1(new_n1102), .A2(new_n1104), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n1118), .B2(new_n537), .ZN(new_n1119));
  AOI211_X1 g694(.A(KEYINPUT59), .B(new_n536), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1112), .A2(new_n1098), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1087), .A2(KEYINPUT124), .A3(new_n1097), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT124), .B1(new_n1087), .B2(new_n1097), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1099), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(new_n799), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n799), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1108), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1111), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G168), .A2(new_n1062), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1075), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1135), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n687), .A2(new_n1063), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT51), .B(new_n1137), .C1(new_n1138), .C2(new_n1062), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  NOR4_X1   g715(.A1(new_n1138), .A2(new_n1140), .A3(new_n1062), .A4(G168), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT125), .B1(new_n1075), .B2(G286), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1136), .B(new_n1139), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n1035), .B2(new_n737), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n726), .B2(new_n1033), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n469), .B(KEYINPUT126), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n470), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n737), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1148));
  NOR4_X1   g723(.A1(new_n987), .A2(new_n467), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1069), .ZN(new_n1150));
  XNOR2_X1  g725(.A(G171), .B(KEYINPUT54), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1145), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n737), .A2(KEYINPUT53), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1072), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1145), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1061), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1082), .B1(new_n1133), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1145), .A2(new_n1154), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1061), .A2(new_n1159), .A3(G301), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1143), .B2(KEYINPUT62), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1075), .A2(G286), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1140), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1075), .A2(KEYINPUT125), .A3(G286), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1162), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1005), .B1(new_n1158), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n990), .B1(new_n996), .B2(new_n696), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT46), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(new_n995), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1172), .B2(new_n995), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT47), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n998), .A2(new_n1001), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n813), .A2(new_n1106), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n990), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n990), .A2(G290), .A3(G1986), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT48), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1003), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1175), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1170), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g758(.A(G319), .ZN(new_n1185));
  NOR4_X1   g759(.A1(G229), .A2(G227), .A3(new_n1185), .A4(G401), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n965), .A2(new_n885), .A3(new_n1186), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


