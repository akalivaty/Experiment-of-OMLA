//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT69), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n468), .B(new_n473), .C1(new_n470), .C2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(new_n469), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n470), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n472), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n479), .A2(KEYINPUT70), .A3(G124), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n482), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(G162));
  NAND2_X1  g063(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n470), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n466), .A2(G102), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n489), .A2(new_n491), .A3(G138), .A4(new_n470), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n469), .A2(G138), .A3(new_n470), .A4(new_n502), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(G62), .A3(G651), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n512), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n509), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n523), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NOR2_X1   g103(.A1(new_n519), .A2(new_n509), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n512), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n529), .A2(G52), .B1(G651), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n520), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n512), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n520), .A2(G81), .B1(G651), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT75), .B(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n529), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT77), .ZN(G188));
  AOI22_X1  g134(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n515), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n520), .B2(G91), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n524), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n529), .A2(KEYINPUT9), .A3(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT78), .B1(new_n566), .B2(new_n567), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n529), .A2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n520), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n524), .A2(G86), .A3(new_n513), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n520), .A2(new_n579), .A3(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n512), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n529), .A2(G48), .B1(G651), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n520), .A2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n529), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n587), .B(new_n588), .C1(new_n515), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n521), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n512), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n529), .A2(G54), .B1(G651), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT10), .B1(new_n521), .B2(new_n592), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  XOR2_X1   g178(.A(G299), .B(KEYINPUT80), .Z(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n469), .A2(new_n466), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  NOR2_X1   g190(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  OR3_X1    g193(.A1(new_n480), .A2(KEYINPUT82), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n472), .A2(G135), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT82), .B1(new_n480), .B2(new_n618), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n619), .A2(new_n620), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n624), .A2(G2096), .B1(KEYINPUT81), .B2(G2100), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n617), .B(new_n625), .C1(G2096), .C2(new_n624), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT17), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  INV_X1    g225(.A(new_n641), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(KEYINPUT84), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(KEYINPUT84), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n649), .B(new_n650), .C1(new_n646), .C2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(G227));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  AOI22_X1  g245(.A1(new_n668), .A2(new_n669), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n665), .A2(new_n670), .A3(new_n667), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n671), .B(new_n672), .C1(new_n669), .C2(new_n668), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT22), .B(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  AND2_X1   g254(.A1(KEYINPUT87), .A2(G29), .ZN(new_n680));
  NOR2_X1   g255(.A1(KEYINPUT87), .A2(G29), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G26), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT92), .Z(new_n685));
  OR2_X1    g260(.A1(new_n685), .A2(KEYINPUT28), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(KEYINPUT28), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n479), .A2(G128), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n472), .A2(G140), .ZN(new_n690));
  OR2_X1    g265(.A1(G104), .A2(G2105), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n691), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n686), .B(new_n687), .C1(new_n688), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2067), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n701), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT34), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n683), .A2(G25), .ZN(new_n712));
  NOR2_X1   g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT88), .Z(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n472), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n479), .A2(G119), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n712), .B1(new_n719), .B2(new_n683), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT89), .B(G1986), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n711), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n726), .A2(new_n728), .ZN(new_n731));
  NAND2_X1  g306(.A1(G168), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G16), .B2(G21), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT95), .B(G1966), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2072), .ZN(new_n737));
  OR2_X1    g312(.A1(G29), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n466), .A2(G103), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT25), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n472), .A2(G139), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n741), .B(new_n742), .C1(new_n470), .C2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n688), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n736), .B1(new_n737), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT24), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(G34), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(G34), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n683), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n475), .B2(new_n688), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n746), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n698), .A2(G20), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT98), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT23), .ZN(new_n756));
  INV_X1    g331(.A(G299), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n698), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n698), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n551), .B2(new_n698), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1341), .Z(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n479), .A2(G129), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n472), .A2(G141), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n466), .A2(G105), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n753), .A2(new_n760), .A3(new_n763), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G4), .B2(G16), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n778), .A2(G4), .A3(G16), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n779), .B(new_n780), .C1(new_n599), .C2(new_n698), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1348), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n683), .A2(G27), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n683), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n745), .A2(new_n737), .B1(G2078), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n785), .C1(G2078), .C2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n698), .A2(G5), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G171), .B2(new_n698), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT97), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n733), .A2(new_n735), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n688), .B1(new_n793), .B2(G28), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(G28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n792), .B(new_n799), .C1(new_n747), .C2(new_n752), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n786), .A2(new_n791), .A3(new_n800), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n730), .A2(new_n731), .A3(new_n777), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n624), .A2(new_n683), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n682), .A2(G35), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n682), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT29), .B(G2090), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n697), .A2(new_n802), .A3(new_n804), .A4(new_n808), .ZN(G311));
  NAND4_X1  g384(.A1(new_n802), .A2(new_n697), .A3(new_n804), .A4(new_n808), .ZN(G150));
  NAND2_X1  g385(.A1(new_n520), .A2(G93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n529), .A2(G55), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n811), .B(new_n812), .C1(new_n515), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT99), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n551), .B(new_n814), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n599), .A2(new_n607), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n817), .B1(new_n822), .B2(G860), .ZN(G145));
  OAI21_X1  g398(.A(KEYINPUT101), .B1(new_n494), .B2(new_n496), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n469), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n495), .C1(new_n826), .C2(new_n470), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT100), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT100), .B1(new_n504), .B2(new_n505), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n824), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n693), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n771), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(KEYINPUT102), .B2(new_n744), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n744), .B(KEYINPUT102), .Z(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n833), .ZN(new_n836));
  INV_X1    g411(.A(G142), .ZN(new_n837));
  NOR2_X1   g412(.A1(G106), .A2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n471), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G130), .B2(new_n479), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n614), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n718), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n836), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(G160), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n624), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g425(.A1(G299), .A2(new_n600), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n562), .B(new_n599), .C1(new_n570), .C2(new_n571), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(G299), .A2(KEYINPUT103), .A3(new_n600), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n851), .A2(new_n853), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT41), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(KEYINPUT41), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n609), .B(new_n818), .ZN(new_n861));
  MUX2_X1   g436(.A(new_n856), .B(new_n860), .S(new_n861), .Z(new_n862));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n865));
  XNOR2_X1  g440(.A(G290), .B(KEYINPUT104), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G305), .ZN(new_n867));
  XNOR2_X1  g442(.A(G303), .B(G288), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n864), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n862), .B(KEYINPUT42), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(KEYINPUT105), .A3(new_n869), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n873), .A3(G868), .ZN(new_n874));
  INV_X1    g449(.A(G868), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT106), .B1(new_n814), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT106), .A4(G868), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(G295));
  AND2_X1   g454(.A1(new_n877), .A2(new_n878), .ZN(G331));
  XOR2_X1   g455(.A(G286), .B(G301), .Z(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n818), .Z(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n858), .B2(new_n859), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n881), .B(new_n818), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n855), .B2(new_n854), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n883), .A2(KEYINPUT107), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT107), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n869), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n848), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT108), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n870), .B1(new_n883), .B2(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n892), .A3(new_n848), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n890), .A2(KEYINPUT43), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n884), .A2(KEYINPUT41), .B1(new_n855), .B2(new_n854), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n884), .A2(KEYINPUT41), .A3(new_n857), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n869), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n891), .B(new_n848), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n899), .A2(new_n900), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n900), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n905), .B2(new_n895), .ZN(G397));
  INV_X1    g481(.A(G1384), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT45), .B1(new_n830), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G40), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n475), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(G1996), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n771), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n911), .B(KEYINPUT109), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G2067), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n693), .B(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(G1996), .B2(new_n770), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n913), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n718), .B(new_n721), .Z(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(G290), .B(G1986), .Z(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n911), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n830), .A2(new_n925), .A3(new_n907), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n830), .B2(new_n907), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n910), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G8), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n706), .A2(G1976), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT52), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(KEYINPUT113), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1976), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT52), .B1(G288), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT114), .Z(new_n939));
  AND2_X1   g514(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n939), .A2(new_n932), .A3(new_n933), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1981), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n581), .A2(new_n943), .A3(new_n585), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n585), .A2(new_n577), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(G1981), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n944), .A2(KEYINPUT49), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT49), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n936), .A2(new_n942), .B1(new_n932), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G8), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT55), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n507), .A2(new_n907), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n830), .A2(new_n907), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n955), .B(new_n910), .C1(new_n956), .C2(new_n954), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(G1971), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(KEYINPUT111), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n830), .A2(new_n925), .A3(new_n907), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n929), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n953), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n497), .B2(new_n506), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n964), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(G2090), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n952), .B(G8), .C1(new_n960), .C2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n960), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n964), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n910), .C1(new_n963), .C2(new_n964), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n978), .A2(G2090), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n931), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n950), .B(new_n973), .C1(new_n952), .C2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n965), .A2(new_n983), .A3(new_n747), .A4(new_n970), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n964), .B1(new_n926), .B2(new_n927), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n985), .A2(new_n747), .A3(new_n910), .A4(new_n970), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT117), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n910), .B1(new_n954), .B2(new_n953), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n734), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n984), .A2(new_n987), .A3(G168), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n931), .A2(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT51), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G8), .A3(G286), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n997), .A3(new_n992), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g575(.A(G2078), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT53), .B1(new_n959), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n790), .B2(new_n971), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n988), .A2(new_n989), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1001), .A2(KEYINPUT53), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT62), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n994), .A2(new_n1008), .A3(new_n996), .A4(new_n998), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1000), .A2(G171), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(G301), .B(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n910), .B1(new_n956), .B2(new_n954), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(new_n908), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1012), .B1(new_n1015), .B2(new_n1005), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1003), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n999), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n562), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n568), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT56), .B(G2072), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n957), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n978), .B2(new_n759), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(KEYINPUT118), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(new_n1026), .C1(new_n978), .C2(new_n759), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1023), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1348), .B1(new_n965), .B2(new_n970), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n930), .A2(new_n916), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n599), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT119), .B(new_n1023), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1033), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1027), .A2(new_n1022), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1041), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT61), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1027), .B2(new_n1022), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1043), .B(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT121), .B(G1341), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT58), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n928), .B2(new_n929), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT120), .B(G1996), .Z(new_n1050));
  OR2_X1    g625(.A1(new_n957), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n551), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1036), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1058), .A2(new_n1034), .A3(KEYINPUT60), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1056), .A2(new_n1057), .B1(new_n1059), .B2(new_n600), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1058), .A2(new_n1034), .A3(new_n600), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT60), .B1(new_n1037), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1057), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1063), .A2(new_n551), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1046), .A2(new_n1060), .A3(new_n1062), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1018), .B1(new_n1042), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n982), .B1(new_n1011), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n995), .A2(G8), .A3(G168), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n981), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n972), .B2(new_n960), .ZN(new_n1073));
  INV_X1    g648(.A(new_n952), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1071), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n973), .A3(new_n950), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n949), .A2(new_n932), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n937), .A3(new_n706), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n944), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n932), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n936), .A2(new_n942), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1084), .B2(new_n973), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT115), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1087), .C1(new_n1084), .C2(new_n973), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1078), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n924), .B1(new_n1069), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(new_n912), .B(KEYINPUT46), .Z(new_n1092));
  OAI21_X1  g667(.A(new_n914), .B1(new_n770), .B2(new_n918), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT47), .Z(new_n1095));
  INV_X1    g670(.A(new_n920), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n721), .A3(new_n719), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n693), .A2(G2067), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n915), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n911), .A2(G1986), .A3(G290), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n1101), .B(KEYINPUT48), .Z(new_n1102));
  AND2_X1   g677(.A1(new_n922), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1095), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT125), .B1(new_n1091), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1078), .A2(new_n1089), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1060), .A2(new_n1066), .A3(new_n1062), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1109), .A2(new_n1046), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1010), .B1(new_n1110), .B2(new_n1018), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1111), .B2(new_n982), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1107), .B(new_n1104), .C1(new_n1112), .C2(new_n924), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1106), .A2(new_n1113), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g689(.A1(G227), .A2(new_n463), .ZN(new_n1116));
  XOR2_X1   g690(.A(new_n1116), .B(KEYINPUT126), .Z(new_n1117));
  NAND2_X1  g691(.A1(new_n1117), .A2(new_n639), .ZN(new_n1118));
  NAND2_X1  g692(.A1(new_n1118), .A2(KEYINPUT127), .ZN(new_n1119));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n1120));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1120), .A3(new_n639), .ZN(new_n1121));
  AOI21_X1  g695(.A(G229), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g696(.A1(new_n1122), .A2(new_n849), .A3(new_n901), .A4(new_n894), .ZN(G225));
  INV_X1    g697(.A(G225), .ZN(G308));
endmodule


