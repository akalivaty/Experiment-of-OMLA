

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n528), .A2(G2104), .ZN(n883) );
  XNOR2_X1 U555 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U556 ( .A1(n705), .A2(n704), .ZN(n708) );
  AND2_X1 U557 ( .A1(n730), .A2(n729), .ZN(n731) );
  INV_X1 U558 ( .A(KEYINPUT17), .ZN(n523) );
  XNOR2_X1 U559 ( .A(n534), .B(n533), .ZN(G164) );
  OR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n520) );
  NOR2_X1 U561 ( .A1(n746), .A2(n804), .ZN(n521) );
  INV_X1 U562 ( .A(n693), .ZN(n723) );
  XNOR2_X1 U563 ( .A(n706), .B(KEYINPUT93), .ZN(n707) );
  XNOR2_X1 U564 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n718) );
  XNOR2_X1 U565 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U566 ( .A1(G8), .A2(n723), .ZN(n804) );
  INV_X1 U567 ( .A(KEYINPUT97), .ZN(n740) );
  NAND2_X1 U568 ( .A1(n880), .A2(G138), .ZN(n525) );
  NOR2_X1 U569 ( .A1(n648), .A2(G651), .ZN(n643) );
  AND2_X1 U570 ( .A1(n820), .A2(n819), .ZN(n821) );
  INV_X1 U571 ( .A(KEYINPUT85), .ZN(n533) );
  NOR2_X1 U572 ( .A1(n532), .A2(n531), .ZN(n534) );
  INV_X1 U573 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U574 ( .A1(n883), .A2(G102), .ZN(n522) );
  XOR2_X1 U575 ( .A(KEYINPUT83), .B(n522), .Z(n526) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XNOR2_X2 U577 ( .A(n524), .B(n523), .ZN(n880) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U579 ( .A(n527), .B(KEYINPUT84), .ZN(n532) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U581 ( .A1(G114), .A2(n875), .ZN(n530) );
  NOR2_X1 U582 ( .A1(G2104), .A2(n528), .ZN(n876) );
  NAND2_X1 U583 ( .A1(G126), .A2(n876), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G113), .A2(n875), .ZN(n536) );
  NAND2_X1 U586 ( .A1(G137), .A2(n880), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U588 ( .A(n537), .B(KEYINPUT65), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G125), .A2(n876), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G101), .A2(n883), .ZN(n540) );
  XNOR2_X1 U592 ( .A(KEYINPUT23), .B(n540), .ZN(n541) );
  NOR2_X1 U593 ( .A1(n542), .A2(n541), .ZN(G160) );
  INV_X1 U594 ( .A(G651), .ZN(n546) );
  NOR2_X1 U595 ( .A1(G543), .A2(n546), .ZN(n543) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n543), .Z(n647) );
  NAND2_X1 U597 ( .A1(G65), .A2(n647), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n648) );
  NAND2_X1 U599 ( .A1(G53), .A2(n643), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n550) );
  NOR2_X1 U601 ( .A1(n648), .A2(n546), .ZN(n633) );
  NAND2_X1 U602 ( .A1(G78), .A2(n633), .ZN(n548) );
  NOR2_X1 U603 ( .A1(G543), .A2(G651), .ZN(n636) );
  NAND2_X1 U604 ( .A1(G91), .A2(n636), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(G299) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U608 ( .A1(n883), .A2(G99), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G111), .A2(n875), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G135), .A2(n880), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n876), .A2(G123), .ZN(n553) );
  XOR2_X1 U613 ( .A(KEYINPUT18), .B(n553), .Z(n554) );
  NOR2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT73), .B(n558), .Z(n924) );
  XNOR2_X1 U617 ( .A(G2096), .B(n924), .ZN(n559) );
  OR2_X1 U618 ( .A1(G2100), .A2(n559), .ZN(G156) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G108), .ZN(G238) );
  NAND2_X1 U622 ( .A1(G75), .A2(n633), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n560), .B(KEYINPUT76), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n647), .A2(G62), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G88), .A2(n636), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G50), .A2(n643), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U629 ( .A1(n566), .A2(n565), .ZN(G166) );
  NAND2_X1 U630 ( .A1(G64), .A2(n647), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G52), .A2(n643), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G77), .A2(n633), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G90), .A2(n636), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(G171) );
  NAND2_X1 U638 ( .A1(n636), .A2(G89), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G76), .A2(n633), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT5), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G63), .A2(n647), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G51), .A2(n643), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT6), .B(n580), .Z(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U652 ( .A(G223), .ZN(n822) );
  NAND2_X1 U653 ( .A1(n822), .A2(G567), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U655 ( .A1(G56), .A2(n647), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n586), .Z(n592) );
  NAND2_X1 U657 ( .A1(n636), .A2(G81), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G68), .A2(n633), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n643), .A2(G43), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n988) );
  INV_X1 U665 ( .A(G860), .ZN(n609) );
  OR2_X1 U666 ( .A1(n988), .A2(n609), .ZN(G153) );
  INV_X1 U667 ( .A(G171), .ZN(G301) );
  INV_X1 U668 ( .A(G868), .ZN(n660) );
  NOR2_X1 U669 ( .A1(G301), .A2(n660), .ZN(n605) );
  NAND2_X1 U670 ( .A1(G54), .A2(n643), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G79), .A2(n633), .ZN(n596) );
  NAND2_X1 U672 ( .A1(G66), .A2(n647), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G92), .A2(n636), .ZN(n597) );
  XNOR2_X1 U675 ( .A(KEYINPUT69), .B(n597), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT15), .ZN(n603) );
  XOR2_X1 U679 ( .A(KEYINPUT70), .B(n603), .Z(n972) );
  NOR2_X1 U680 ( .A1(n972), .A2(G868), .ZN(n604) );
  NOR2_X1 U681 ( .A1(n605), .A2(n604), .ZN(G284) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT71), .B(n606), .Z(n608) );
  NOR2_X1 U684 ( .A1(G286), .A2(n660), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U686 ( .A1(G559), .A2(n609), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT72), .ZN(n611) );
  INV_X1 U688 ( .A(n972), .ZN(n898) );
  NAND2_X1 U689 ( .A1(n611), .A2(n898), .ZN(n612) );
  XNOR2_X1 U690 ( .A(KEYINPUT16), .B(n612), .ZN(G148) );
  NOR2_X1 U691 ( .A1(G868), .A2(n988), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n898), .A2(G868), .ZN(n613) );
  NOR2_X1 U693 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U694 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G67), .A2(n647), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G93), .A2(n636), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G80), .A2(n633), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G55), .A2(n643), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n659) );
  NAND2_X1 U702 ( .A1(n898), .A2(G559), .ZN(n622) );
  XOR2_X1 U703 ( .A(n988), .B(n622), .Z(n657) );
  XOR2_X1 U704 ( .A(n657), .B(KEYINPUT74), .Z(n623) );
  NOR2_X1 U705 ( .A1(G860), .A2(n623), .ZN(n624) );
  XOR2_X1 U706 ( .A(KEYINPUT75), .B(n624), .Z(n625) );
  XOR2_X1 U707 ( .A(n659), .B(n625), .Z(G145) );
  NAND2_X1 U708 ( .A1(G61), .A2(n647), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G86), .A2(n636), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n633), .A2(G73), .ZN(n628) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(n628), .Z(n629) );
  NOR2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n643), .A2(G48), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U716 ( .A1(n643), .A2(G47), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G72), .A2(n633), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G60), .A2(n647), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n636), .A2(G85), .ZN(n637) );
  XOR2_X1 U721 ( .A(KEYINPUT66), .B(n637), .Z(n638) );
  NOR2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U724 ( .A(KEYINPUT67), .B(n642), .Z(G290) );
  NAND2_X1 U725 ( .A1(G49), .A2(n643), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(G288) );
  XOR2_X1 U731 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n651) );
  XNOR2_X1 U732 ( .A(G299), .B(n651), .ZN(n654) );
  XNOR2_X1 U733 ( .A(G166), .B(G305), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n652), .B(G290), .ZN(n653) );
  XNOR2_X1 U735 ( .A(n654), .B(n653), .ZN(n656) );
  XOR2_X1 U736 ( .A(G288), .B(n659), .Z(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n895) );
  XNOR2_X1 U738 ( .A(n657), .B(n895), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n664), .ZN(n666) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(KEYINPUT78), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U747 ( .A1(G2072), .A2(n667), .ZN(G158) );
  XOR2_X1 U748 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n668) );
  NOR2_X1 U752 ( .A1(G237), .A2(n668), .ZN(n669) );
  XOR2_X1 U753 ( .A(KEYINPUT80), .B(n669), .Z(n670) );
  NOR2_X1 U754 ( .A1(G238), .A2(n670), .ZN(n671) );
  XNOR2_X1 U755 ( .A(KEYINPUT81), .B(n671), .ZN(n828) );
  NAND2_X1 U756 ( .A1(G567), .A2(n828), .ZN(n677) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n672) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U759 ( .A1(G218), .A2(n673), .ZN(n674) );
  XOR2_X1 U760 ( .A(KEYINPUT79), .B(n674), .Z(n675) );
  NAND2_X1 U761 ( .A1(G96), .A2(n675), .ZN(n827) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n827), .ZN(n676) );
  NAND2_X1 U763 ( .A1(n677), .A2(n676), .ZN(n849) );
  NOR2_X1 U764 ( .A1(n678), .A2(n849), .ZN(n679) );
  XNOR2_X1 U765 ( .A(n679), .B(KEYINPUT82), .ZN(n825) );
  NAND2_X1 U766 ( .A1(G36), .A2(n825), .ZN(G176) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n769) );
  NOR2_X1 U769 ( .A1(n520), .A2(n769), .ZN(n680) );
  XNOR2_X1 U770 ( .A(n680), .B(KEYINPUT64), .ZN(n693) );
  XOR2_X1 U771 ( .A(G2078), .B(KEYINPUT25), .Z(n681) );
  XNOR2_X1 U772 ( .A(KEYINPUT90), .B(n681), .ZN(n955) );
  NAND2_X1 U773 ( .A1(n693), .A2(n955), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n723), .A2(G1961), .ZN(n682) );
  NAND2_X1 U775 ( .A1(n683), .A2(n682), .ZN(n714) );
  OR2_X1 U776 ( .A1(n714), .A2(G301), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n723), .A2(G1348), .ZN(n685) );
  NAND2_X1 U778 ( .A1(G2067), .A2(n693), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U780 ( .A(n686), .B(KEYINPUT92), .Z(n692) );
  AND2_X1 U781 ( .A1(n898), .A2(n692), .ZN(n691) );
  NAND2_X1 U782 ( .A1(G2072), .A2(n693), .ZN(n687) );
  XOR2_X1 U783 ( .A(KEYINPUT27), .B(n687), .Z(n689) );
  XOR2_X1 U784 ( .A(G1956), .B(KEYINPUT91), .Z(n1002) );
  NAND2_X1 U785 ( .A1(n723), .A2(n1002), .ZN(n688) );
  NAND2_X1 U786 ( .A1(n689), .A2(n688), .ZN(n702) );
  NOR2_X1 U787 ( .A1(n702), .A2(G299), .ZN(n690) );
  NOR2_X1 U788 ( .A1(n691), .A2(n690), .ZN(n701) );
  OR2_X1 U789 ( .A1(n898), .A2(n692), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n693), .A2(G1996), .ZN(n694) );
  XNOR2_X1 U791 ( .A(n694), .B(KEYINPUT26), .ZN(n696) );
  NAND2_X1 U792 ( .A1(n723), .A2(G1341), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n988), .A2(n697), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n705) );
  AND2_X1 U797 ( .A1(G299), .A2(n702), .ZN(n703) );
  XNOR2_X1 U798 ( .A(KEYINPUT28), .B(n703), .ZN(n704) );
  INV_X1 U799 ( .A(KEYINPUT29), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n721) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n804), .ZN(n735) );
  NOR2_X1 U802 ( .A1(n723), .A2(G2084), .ZN(n732) );
  NOR2_X1 U803 ( .A1(n735), .A2(n732), .ZN(n711) );
  NAND2_X1 U804 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U805 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U806 ( .A1(G168), .A2(n713), .ZN(n717) );
  NAND2_X1 U807 ( .A1(G301), .A2(n714), .ZN(n715) );
  XOR2_X1 U808 ( .A(KEYINPUT94), .B(n715), .Z(n716) );
  NOR2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n733) );
  NAND2_X1 U811 ( .A1(n733), .A2(G286), .ZN(n730) );
  INV_X1 U812 ( .A(G8), .ZN(n728) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n804), .ZN(n722) );
  XNOR2_X1 U814 ( .A(n722), .B(KEYINPUT96), .ZN(n725) );
  NOR2_X1 U815 ( .A1(n723), .A2(G2090), .ZN(n724) );
  NOR2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G303), .A2(n726), .ZN(n727) );
  OR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n731), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U820 ( .A1(G8), .A2(n732), .ZN(n737) );
  INV_X1 U821 ( .A(n733), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U825 ( .A(n741), .B(n740), .ZN(n802) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U828 ( .A1(n975), .A2(n742), .ZN(n744) );
  INV_X1 U829 ( .A(KEYINPUT33), .ZN(n743) );
  AND2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n802), .A2(n745), .ZN(n775) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n976) );
  INV_X1 U833 ( .A(n976), .ZN(n746) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n521), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n975), .A2(KEYINPUT33), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n804), .A2(n747), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n773) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n969) );
  NAND2_X1 U839 ( .A1(G119), .A2(n876), .ZN(n751) );
  NAND2_X1 U840 ( .A1(G95), .A2(n883), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n880), .A2(G131), .ZN(n752) );
  XOR2_X1 U843 ( .A(KEYINPUT86), .B(n752), .Z(n753) );
  NOR2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n875), .A2(G107), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n887) );
  NAND2_X1 U847 ( .A1(G1991), .A2(n887), .ZN(n757) );
  XNOR2_X1 U848 ( .A(n757), .B(KEYINPUT87), .ZN(n768) );
  NAND2_X1 U849 ( .A1(G105), .A2(n883), .ZN(n758) );
  XNOR2_X1 U850 ( .A(n758), .B(KEYINPUT38), .ZN(n763) );
  NAND2_X1 U851 ( .A1(G117), .A2(n875), .ZN(n760) );
  NAND2_X1 U852 ( .A1(G129), .A2(n876), .ZN(n759) );
  NAND2_X1 U853 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U854 ( .A(KEYINPUT88), .B(n761), .Z(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U856 ( .A1(G141), .A2(n880), .ZN(n764) );
  XNOR2_X1 U857 ( .A(KEYINPUT89), .B(n764), .ZN(n765) );
  OR2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n874) );
  AND2_X1 U859 ( .A1(G1996), .A2(n874), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n776) );
  XOR2_X1 U861 ( .A(G1986), .B(G290), .Z(n981) );
  NAND2_X1 U862 ( .A1(n776), .A2(n981), .ZN(n771) );
  INV_X1 U863 ( .A(n520), .ZN(n770) );
  NOR2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n816) );
  NAND2_X1 U865 ( .A1(n771), .A2(n816), .ZN(n807) );
  AND2_X1 U866 ( .A1(n969), .A2(n807), .ZN(n772) );
  AND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n796) );
  NOR2_X1 U869 ( .A1(G1996), .A2(n874), .ZN(n929) );
  INV_X1 U870 ( .A(n776), .ZN(n921) );
  NOR2_X1 U871 ( .A1(n887), .A2(G1991), .ZN(n777) );
  XNOR2_X1 U872 ( .A(n777), .B(KEYINPUT98), .ZN(n927) );
  NOR2_X1 U873 ( .A1(G1986), .A2(G290), .ZN(n778) );
  NOR2_X1 U874 ( .A1(n927), .A2(n778), .ZN(n779) );
  NOR2_X1 U875 ( .A1(n921), .A2(n779), .ZN(n780) );
  NOR2_X1 U876 ( .A1(n929), .A2(n780), .ZN(n781) );
  XOR2_X1 U877 ( .A(n781), .B(KEYINPUT39), .Z(n782) );
  XNOR2_X1 U878 ( .A(KEYINPUT99), .B(n782), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n783), .A2(n816), .ZN(n794) );
  XOR2_X1 U880 ( .A(G2067), .B(KEYINPUT37), .Z(n815) );
  NAND2_X1 U881 ( .A1(G140), .A2(n880), .ZN(n785) );
  NAND2_X1 U882 ( .A1(G104), .A2(n883), .ZN(n784) );
  NAND2_X1 U883 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U885 ( .A1(G116), .A2(n875), .ZN(n788) );
  NAND2_X1 U886 ( .A1(G128), .A2(n876), .ZN(n787) );
  NAND2_X1 U887 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U888 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U889 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U890 ( .A(KEYINPUT36), .B(n792), .Z(n892) );
  NOR2_X1 U891 ( .A1(n815), .A2(n892), .ZN(n793) );
  XNOR2_X1 U892 ( .A(n793), .B(KEYINPUT100), .ZN(n943) );
  NAND2_X1 U893 ( .A1(n943), .A2(n816), .ZN(n814) );
  AND2_X1 U894 ( .A1(n794), .A2(n814), .ZN(n795) );
  AND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n813) );
  NAND2_X1 U896 ( .A1(G8), .A2(G166), .ZN(n797) );
  NOR2_X1 U897 ( .A1(G2090), .A2(n797), .ZN(n800) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XOR2_X1 U899 ( .A(n798), .B(KEYINPUT24), .Z(n799) );
  NOR2_X1 U900 ( .A1(n804), .A2(n799), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n800), .A2(n803), .ZN(n801) );
  NAND2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n811) );
  INV_X1 U903 ( .A(n803), .ZN(n806) );
  INV_X1 U904 ( .A(n804), .ZN(n805) );
  AND2_X1 U905 ( .A1(n806), .A2(n805), .ZN(n809) );
  INV_X1 U906 ( .A(n807), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n820) );
  INV_X1 U910 ( .A(n814), .ZN(n818) );
  AND2_X1 U911 ( .A1(n892), .A2(n815), .ZN(n922) );
  NAND2_X1 U912 ( .A1(n922), .A2(n816), .ZN(n817) );
  OR2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U914 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U917 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT104), .B(n826), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(G2474), .B(G1981), .Z(n830) );
  XNOR2_X1 U928 ( .A(G1966), .B(G1961), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U930 ( .A(n831), .B(KEYINPUT107), .Z(n833) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U933 ( .A(G1986), .B(G1976), .Z(n835) );
  XNOR2_X1 U934 ( .A(G1956), .B(G1971), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U936 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2072), .B(G2678), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n842), .B(KEYINPUT42), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT106), .B(G2100), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(G227) );
  INV_X1 U949 ( .A(n849), .ZN(G319) );
  NAND2_X1 U950 ( .A1(G124), .A2(n876), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n875), .A2(G112), .ZN(n851) );
  NAND2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G136), .A2(n880), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G100), .A2(n883), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U957 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G118), .A2(n875), .ZN(n865) );
  NAND2_X1 U959 ( .A1(n876), .A2(G130), .ZN(n857) );
  XNOR2_X1 U960 ( .A(KEYINPUT109), .B(n857), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G142), .A2(n880), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G106), .A2(n883), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U964 ( .A(KEYINPUT45), .B(n860), .Z(n861) );
  XNOR2_X1 U965 ( .A(KEYINPUT110), .B(n861), .ZN(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n867) );
  XNOR2_X1 U969 ( .A(G162), .B(KEYINPUT46), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT113), .B(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n924), .B(KEYINPUT114), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n891) );
  NAND2_X1 U976 ( .A1(G115), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G127), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n879), .B(KEYINPUT47), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U982 ( .A1(G103), .A2(n883), .ZN(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT111), .B(n884), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n934) );
  XNOR2_X1 U985 ( .A(n887), .B(n934), .ZN(n889) );
  XNOR2_X1 U986 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U990 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n895), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n988), .B(G171), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n900) );
  XOR2_X1 U994 ( .A(n898), .B(KEYINPUT115), .Z(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n903) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n917) );
  XOR2_X1 U1000 ( .A(KEYINPUT103), .B(G2446), .Z(n905) );
  XNOR2_X1 U1001 ( .A(KEYINPUT101), .B(G2451), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n906), .B(G2430), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1006 ( .A(KEYINPUT102), .B(G2438), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G2435), .B(G2454), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2427), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n915), .A2(G14), .ZN(n920) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n920), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n941) );
  XOR2_X1 U1020 ( .A(G160), .B(G2084), .Z(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT117), .B(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT118), .B(n928), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n931), .Z(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n939) );
  XOR2_X1 U1029 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n937), .Z(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n965) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n965), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(G29), .ZN(n1029) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n960) );
  XNOR2_X1 U1041 ( .A(G2072), .B(G33), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1991), .B(G25), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n949) );
  NAND2_X1 U1045 ( .A1(n949), .A2(G28), .ZN(n952) );
  XOR2_X1 U1046 ( .A(G32), .B(G1996), .Z(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT119), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G27), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n967) );
  INV_X1 U1058 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n968), .ZN(n1027) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(KEYINPUT57), .ZN(n993) );
  XNOR2_X1 U1065 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n972), .B(G1348), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n987) );
  INV_X1 U1068 ( .A(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G299), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G1971), .B(KEYINPUT120), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n982), .B(G303), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT121), .B(n985), .Z(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n988), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT122), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n1025) );
  INV_X1 U1083 ( .A(G16), .ZN(n1023) );
  XOR2_X1 U1084 ( .A(G1986), .B(G24), .Z(n999) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G22), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(G23), .B(G1976), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(n1001), .B(n1000), .ZN(n1020) );
  XOR2_X1 U1091 ( .A(G1961), .B(G5), .Z(n1015) );
  XNOR2_X1 U1092 ( .A(n1002), .B(G20), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT123), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT124), .B(n1008), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G1348), .B(KEYINPUT59), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(G4), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(n1012), .B(KEYINPUT125), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT60), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT126), .B(G1966), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(G21), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1021), .Z(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

