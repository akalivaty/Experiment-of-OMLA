

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768;

  AND2_X1 U373 ( .A1(n598), .A2(n349), .ZN(n610) );
  NOR2_X1 U374 ( .A1(n351), .A2(n350), .ZN(n349) );
  AND2_X1 U375 ( .A1(n348), .A2(n596), .ZN(n597) );
  INV_X1 U376 ( .A(n692), .ZN(n350) );
  INV_X1 U377 ( .A(n702), .ZN(n351) );
  XNOR2_X1 U378 ( .A(n404), .B(n403), .ZN(n596) );
  XNOR2_X1 U379 ( .A(n383), .B(n465), .ZN(n731) );
  NOR2_X1 U380 ( .A1(n707), .A2(n565), .ZN(n569) );
  XNOR2_X1 U381 ( .A(n497), .B(n496), .ZN(n501) );
  XNOR2_X1 U382 ( .A(n470), .B(n469), .ZN(n759) );
  XNOR2_X1 U383 ( .A(n472), .B(KEYINPUT10), .ZN(n643) );
  XNOR2_X1 U384 ( .A(G140), .B(G113), .ZN(n502) );
  NOR2_X1 U385 ( .A1(G953), .A2(G237), .ZN(n495) );
  AND2_X2 U386 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X2 U387 ( .A(n378), .B(n533), .ZN(n640) );
  INV_X1 U388 ( .A(n596), .ZN(n728) );
  INV_X1 U389 ( .A(n694), .ZN(n348) );
  XNOR2_X2 U390 ( .A(n507), .B(n508), .ZN(n545) );
  INV_X1 U391 ( .A(G953), .ZN(n473) );
  NAND2_X2 U392 ( .A1(n395), .A2(n392), .ZN(n354) );
  XNOR2_X2 U393 ( .A(G128), .B(G119), .ZN(n432) );
  AND2_X4 U394 ( .A1(n408), .A2(n406), .ZN(n743) );
  AND2_X2 U395 ( .A1(n405), .A2(n409), .ZN(n408) );
  NOR2_X2 U396 ( .A1(n766), .A2(n767), .ZN(n590) );
  NAND2_X1 U397 ( .A1(n407), .A2(KEYINPUT82), .ZN(n406) );
  BUF_X1 U398 ( .A(n640), .Z(n355) );
  AND2_X1 U399 ( .A1(n377), .A2(n373), .ZN(n372) );
  NAND2_X1 U400 ( .A1(n394), .A2(n357), .ZN(n392) );
  NAND2_X2 U401 ( .A1(n390), .A2(n386), .ZN(n580) );
  XNOR2_X1 U402 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U403 ( .A(n661), .B(n660), .ZN(n662) );
  AND2_X1 U404 ( .A1(n381), .A2(n391), .ZN(n390) );
  XNOR2_X1 U405 ( .A(n369), .B(G146), .ZN(n463) );
  NAND2_X1 U406 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U407 ( .A(G128), .B(G143), .ZN(n352) );
  BUF_X1 U408 ( .A(n380), .Z(n353) );
  XNOR2_X1 U409 ( .A(n580), .B(n356), .ZN(n380) );
  NOR2_X2 U410 ( .A1(n553), .A2(KEYINPUT44), .ZN(n526) );
  BUF_X1 U411 ( .A(n535), .Z(n539) );
  INV_X1 U412 ( .A(KEYINPUT84), .ZN(n417) );
  XNOR2_X1 U413 ( .A(G134), .B(G131), .ZN(n458) );
  XNOR2_X1 U414 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n423) );
  INV_X1 U415 ( .A(G140), .ZN(n429) );
  XNOR2_X1 U416 ( .A(G104), .B(G107), .ZN(n425) );
  INV_X1 U417 ( .A(KEYINPUT19), .ZN(n393) );
  NAND2_X1 U418 ( .A1(n599), .A2(KEYINPUT19), .ZN(n396) );
  NOR2_X1 U419 ( .A1(n578), .A2(n579), .ZN(n368) );
  INV_X1 U420 ( .A(KEYINPUT67), .ZN(n375) );
  AND2_X1 U421 ( .A1(n374), .A2(n713), .ZN(n373) );
  NAND2_X1 U422 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U423 ( .A(n530), .ZN(n376) );
  INV_X1 U424 ( .A(KEYINPUT107), .ZN(n403) );
  INV_X1 U425 ( .A(KEYINPUT73), .ZN(n415) );
  INV_X1 U426 ( .A(G237), .ZN(n480) );
  INV_X1 U427 ( .A(G469), .ZN(n389) );
  NAND2_X1 U428 ( .A1(G902), .A2(G469), .ZN(n391) );
  AND2_X1 U429 ( .A1(n617), .A2(n412), .ZN(n411) );
  NOR2_X1 U430 ( .A1(n410), .A2(n703), .ZN(n409) );
  XNOR2_X1 U431 ( .A(G107), .B(G116), .ZN(n511) );
  XNOR2_X1 U432 ( .A(n402), .B(n400), .ZN(n509) );
  XNOR2_X1 U433 ( .A(KEYINPUT78), .B(KEYINPUT8), .ZN(n402) );
  NOR2_X1 U434 ( .A1(n401), .A2(G953), .ZN(n400) );
  INV_X1 U435 ( .A(G234), .ZN(n401) );
  XOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n497) );
  XOR2_X1 U437 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n499) );
  XNOR2_X1 U438 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n475) );
  XNOR2_X1 U439 ( .A(KEYINPUT85), .B(KEYINPUT90), .ZN(n471) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n486) );
  XNOR2_X1 U441 ( .A(G134), .B(G122), .ZN(n514) );
  XOR2_X1 U442 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n515) );
  XNOR2_X1 U443 ( .A(n463), .B(n431), .ZN(n659) );
  XNOR2_X1 U444 ( .A(n586), .B(n585), .ZN(n706) );
  XNOR2_X1 U445 ( .A(n574), .B(n573), .ZN(n618) );
  NAND2_X1 U446 ( .A1(n366), .A2(n572), .ZN(n574) );
  INV_X1 U447 ( .A(KEYINPUT86), .ZN(n379) );
  INV_X1 U448 ( .A(KEYINPUT28), .ZN(n367) );
  XNOR2_X1 U449 ( .A(n716), .B(KEYINPUT6), .ZN(n605) );
  XNOR2_X1 U450 ( .A(n632), .B(KEYINPUT62), .ZN(n633) );
  XNOR2_X1 U451 ( .A(n652), .B(n653), .ZN(n654) );
  XNOR2_X1 U452 ( .A(n636), .B(KEYINPUT87), .ZN(n682) );
  BUF_X1 U453 ( .A(n553), .Z(n673) );
  NAND2_X1 U454 ( .A1(n371), .A2(n375), .ZN(n370) );
  XNOR2_X1 U455 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n356) );
  AND2_X1 U456 ( .A1(n399), .A2(n393), .ZN(n357) );
  AND2_X1 U457 ( .A1(n530), .A2(KEYINPUT67), .ZN(n358) );
  INV_X1 U458 ( .A(G902), .ZN(n388) );
  XNOR2_X2 U459 ( .A(n359), .B(n558), .ZN(n745) );
  NAND2_X1 U460 ( .A1(n362), .A2(n360), .ZN(n359) );
  NOR2_X1 U461 ( .A1(n557), .A2(n361), .ZN(n360) );
  NAND2_X1 U462 ( .A1(n551), .A2(n768), .ZN(n361) );
  XNOR2_X1 U463 ( .A(n363), .B(n415), .ZN(n362) );
  NAND2_X1 U464 ( .A1(n418), .A2(n416), .ZN(n363) );
  NAND2_X1 U465 ( .A1(n640), .A2(n364), .ZN(n552) );
  NAND2_X2 U466 ( .A1(n372), .A2(n370), .ZN(n364) );
  XNOR2_X1 U467 ( .A(n364), .B(G110), .ZN(G12) );
  NOR2_X1 U468 ( .A1(n618), .A2(n696), .ZN(n576) );
  NAND2_X1 U469 ( .A1(n455), .A2(n380), .ZN(n384) );
  NOR2_X2 U470 ( .A1(n384), .A2(n605), .ZN(n383) );
  XNOR2_X2 U471 ( .A(n454), .B(KEYINPUT72), .ZN(n707) );
  XNOR2_X1 U472 ( .A(n369), .B(n478), .ZN(n479) );
  XNOR2_X1 U473 ( .A(n552), .B(n417), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n612), .B(n423), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n365), .B(n435), .ZN(n440) );
  XNOR2_X1 U476 ( .A(n434), .B(n433), .ZN(n365) );
  INV_X1 U477 ( .A(n591), .ZN(n366) );
  NAND2_X1 U478 ( .A1(n569), .A2(n568), .ZN(n591) );
  XNOR2_X1 U479 ( .A(n385), .B(n494), .ZN(n522) );
  XNOR2_X2 U480 ( .A(n441), .B(G902), .ZN(n625) );
  XNOR2_X1 U481 ( .A(n368), .B(n367), .ZN(n582) );
  XNOR2_X2 U482 ( .A(n641), .B(n424), .ZN(n369) );
  INV_X1 U483 ( .A(n414), .ZN(n371) );
  NAND2_X1 U484 ( .A1(n414), .A2(n358), .ZN(n377) );
  NAND2_X1 U485 ( .A1(n414), .A2(n532), .ZN(n378) );
  INV_X1 U486 ( .A(n353), .ZN(n708) );
  XNOR2_X1 U487 ( .A(n708), .B(n379), .ZN(n607) );
  NOR2_X1 U488 ( .A1(n613), .A2(n353), .ZN(n614) );
  NAND2_X1 U489 ( .A1(n659), .A2(G469), .ZN(n381) );
  NAND2_X1 U490 ( .A1(n731), .A2(n382), .ZN(n385) );
  INV_X1 U491 ( .A(n535), .ZN(n382) );
  XNOR2_X2 U492 ( .A(n398), .B(KEYINPUT0), .ZN(n535) );
  XNOR2_X2 U493 ( .A(n510), .B(KEYINPUT4), .ZN(n641) );
  XNOR2_X2 U494 ( .A(G128), .B(G143), .ZN(n510) );
  NOR2_X1 U495 ( .A1(n384), .A2(n579), .ZN(n534) );
  OR2_X1 U496 ( .A1(n659), .A2(n387), .ZN(n386) );
  INV_X1 U497 ( .A(n570), .ZN(n394) );
  NAND2_X1 U498 ( .A1(n570), .A2(KEYINPUT19), .ZN(n397) );
  NAND2_X1 U499 ( .A1(n354), .A2(n493), .ZN(n398) );
  INV_X1 U500 ( .A(n599), .ZN(n399) );
  XNOR2_X2 U501 ( .A(n484), .B(n483), .ZN(n570) );
  NAND2_X1 U502 ( .A1(n619), .A2(n696), .ZN(n404) );
  XNOR2_X1 U503 ( .A(n685), .B(KEYINPUT106), .ZN(n619) );
  XNOR2_X1 U504 ( .A(n543), .B(KEYINPUT105), .ZN(n685) );
  NAND2_X1 U505 ( .A1(n413), .A2(n411), .ZN(n405) );
  INV_X1 U506 ( .A(n413), .ZN(n407) );
  NOR2_X1 U507 ( .A1(n617), .A2(n412), .ZN(n410) );
  INV_X1 U508 ( .A(KEYINPUT82), .ZN(n412) );
  NAND2_X1 U509 ( .A1(n414), .A2(n708), .ZN(n422) );
  XNOR2_X2 U510 ( .A(n529), .B(KEYINPUT22), .ZN(n414) );
  XNOR2_X1 U511 ( .A(n526), .B(n419), .ZN(n418) );
  INV_X1 U512 ( .A(KEYINPUT71), .ZN(n419) );
  XNOR2_X2 U513 ( .A(n421), .B(n420), .ZN(n467) );
  XNOR2_X2 U514 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n420) );
  XNOR2_X2 U515 ( .A(G119), .B(G113), .ZN(n421) );
  XNOR2_X2 U516 ( .A(G146), .B(G125), .ZN(n472) );
  NAND2_X1 U517 ( .A1(n580), .A2(n577), .ZN(n565) );
  XNOR2_X2 U518 ( .A(n631), .B(KEYINPUT65), .ZN(n679) );
  INV_X1 U519 ( .A(n542), .ZN(n544) );
  INV_X1 U520 ( .A(KEYINPUT33), .ZN(n465) );
  INV_X1 U521 ( .A(KEYINPUT74), .ZN(n622) );
  INV_X1 U522 ( .A(n706), .ZN(n739) );
  BUF_X1 U523 ( .A(n666), .Z(n668) );
  XNOR2_X1 U524 ( .A(n525), .B(n524), .ZN(n553) );
  XNOR2_X1 U525 ( .A(KEYINPUT70), .B(G101), .ZN(n424) );
  XNOR2_X1 U526 ( .A(G110), .B(KEYINPUT88), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(n425), .ZN(n428) );
  NAND2_X1 U528 ( .A1(n473), .A2(G227), .ZN(n426) );
  XNOR2_X1 U529 ( .A(n426), .B(KEYINPUT94), .ZN(n427) );
  XNOR2_X1 U530 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U531 ( .A(n429), .B(G137), .ZN(n433) );
  XNOR2_X1 U532 ( .A(n433), .B(n458), .ZN(n642) );
  XNOR2_X1 U533 ( .A(n430), .B(n642), .ZN(n431) );
  NAND2_X1 U534 ( .A1(n509), .A2(G221), .ZN(n435) );
  XNOR2_X1 U535 ( .A(n432), .B(KEYINPUT95), .ZN(n434) );
  XNOR2_X1 U536 ( .A(G110), .B(KEYINPUT23), .ZN(n437) );
  XNOR2_X1 U537 ( .A(KEYINPUT24), .B(KEYINPUT76), .ZN(n436) );
  XNOR2_X1 U538 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U539 ( .A(n643), .B(n438), .ZN(n439) );
  XNOR2_X1 U540 ( .A(n440), .B(n439), .ZN(n675) );
  OR2_X2 U541 ( .A1(n675), .A2(G902), .ZN(n449) );
  INV_X1 U542 ( .A(KEYINPUT15), .ZN(n441) );
  INV_X1 U543 ( .A(n625), .ZN(n442) );
  NAND2_X1 U544 ( .A1(n442), .A2(G234), .ZN(n444) );
  XNOR2_X1 U545 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n443) );
  XNOR2_X1 U546 ( .A(n444), .B(n443), .ZN(n450) );
  AND2_X1 U547 ( .A1(n450), .A2(G217), .ZN(n447) );
  XNOR2_X1 U548 ( .A(KEYINPUT75), .B(KEYINPUT97), .ZN(n445) );
  XNOR2_X1 U549 ( .A(n445), .B(KEYINPUT25), .ZN(n446) );
  XNOR2_X1 U550 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X2 U551 ( .A(n449), .B(n448), .ZN(n548) );
  NAND2_X1 U552 ( .A1(n450), .A2(G221), .ZN(n453) );
  INV_X1 U553 ( .A(KEYINPUT98), .ZN(n451) );
  XNOR2_X1 U554 ( .A(n451), .B(KEYINPUT21), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n453), .B(n452), .ZN(n711) );
  NAND2_X1 U556 ( .A1(n548), .A2(n711), .ZN(n454) );
  INV_X1 U557 ( .A(n707), .ZN(n455) );
  NAND2_X1 U558 ( .A1(n495), .A2(G210), .ZN(n456) );
  XNOR2_X1 U559 ( .A(n456), .B(G137), .ZN(n457) );
  XNOR2_X1 U560 ( .A(n467), .B(n457), .ZN(n461) );
  XOR2_X1 U561 ( .A(G116), .B(KEYINPUT5), .Z(n459) );
  XNOR2_X1 U562 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U563 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n632) );
  OR2_X2 U565 ( .A1(n632), .A2(G902), .ZN(n464) );
  XNOR2_X2 U566 ( .A(n464), .B(G472), .ZN(n716) );
  XNOR2_X2 U567 ( .A(G104), .B(G122), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT16), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n466), .B(n467), .ZN(n470) );
  XNOR2_X1 U570 ( .A(n468), .B(n511), .ZN(n469) );
  XNOR2_X1 U571 ( .A(n472), .B(n471), .ZN(n477) );
  NAND2_X1 U572 ( .A1(n473), .A2(G224), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U574 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U575 ( .A(n479), .B(n759), .ZN(n666) );
  OR2_X2 U576 ( .A1(n666), .A2(n625), .ZN(n484) );
  NAND2_X1 U577 ( .A1(n388), .A2(n480), .ZN(n485) );
  NAND2_X1 U578 ( .A1(n485), .A2(G210), .ZN(n482) );
  INV_X1 U579 ( .A(KEYINPUT91), .ZN(n481) );
  XNOR2_X1 U580 ( .A(n482), .B(n481), .ZN(n483) );
  AND2_X1 U581 ( .A1(n485), .A2(G214), .ZN(n599) );
  XNOR2_X1 U582 ( .A(n486), .B(KEYINPUT92), .ZN(n487) );
  XNOR2_X1 U583 ( .A(KEYINPUT14), .B(n487), .ZN(n491) );
  NAND2_X1 U584 ( .A1(G902), .A2(n491), .ZN(n559) );
  INV_X1 U585 ( .A(n559), .ZN(n490) );
  INV_X1 U586 ( .A(G898), .ZN(n488) );
  NAND2_X1 U587 ( .A1(n488), .A2(G953), .ZN(n489) );
  XNOR2_X1 U588 ( .A(n489), .B(KEYINPUT93), .ZN(n760) );
  NAND2_X1 U589 ( .A1(n490), .A2(n760), .ZN(n492) );
  NAND2_X1 U590 ( .A1(G952), .A2(n491), .ZN(n737) );
  OR2_X1 U591 ( .A1(n737), .A2(G953), .ZN(n562) );
  NAND2_X1 U592 ( .A1(n492), .A2(n562), .ZN(n493) );
  INV_X1 U593 ( .A(KEYINPUT34), .ZN(n494) );
  XNOR2_X1 U594 ( .A(KEYINPUT13), .B(G475), .ZN(n508) );
  NAND2_X1 U595 ( .A1(G214), .A2(n495), .ZN(n496) );
  XNOR2_X1 U596 ( .A(G143), .B(G131), .ZN(n498) );
  XNOR2_X1 U597 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U598 ( .A(n501), .B(n500), .ZN(n506) );
  XNOR2_X1 U599 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U600 ( .A(n643), .B(n504), .ZN(n505) );
  XNOR2_X1 U601 ( .A(n506), .B(n505), .ZN(n652) );
  NOR2_X1 U602 ( .A1(G902), .A2(n652), .ZN(n507) );
  AND2_X1 U603 ( .A1(n509), .A2(G217), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n352), .B(n511), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n519) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT104), .Z(n516) );
  XNOR2_X1 U608 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U609 ( .A(n519), .B(n518), .ZN(n680) );
  NOR2_X1 U610 ( .A1(G902), .A2(n680), .ZN(n520) );
  XNOR2_X2 U611 ( .A(n520), .B(G478), .ZN(n542) );
  AND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n521) );
  XNOR2_X1 U613 ( .A(n521), .B(KEYINPUT110), .ZN(n593) );
  NAND2_X1 U614 ( .A1(n522), .A2(n593), .ZN(n525) );
  INV_X1 U615 ( .A(KEYINPUT77), .ZN(n523) );
  XNOR2_X1 U616 ( .A(n523), .B(KEYINPUT35), .ZN(n524) );
  INV_X1 U617 ( .A(n716), .ZN(n579) );
  AND2_X1 U618 ( .A1(n579), .A2(n708), .ZN(n530) );
  INV_X1 U619 ( .A(n545), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n527), .A2(n542), .ZN(n726) );
  NAND2_X1 U621 ( .A1(n583), .A2(n711), .ZN(n528) );
  NOR2_X2 U622 ( .A1(n535), .A2(n528), .ZN(n529) );
  INV_X1 U623 ( .A(n548), .ZN(n713) );
  AND2_X1 U624 ( .A1(n605), .A2(n713), .ZN(n531) );
  AND2_X1 U625 ( .A1(n607), .A2(n531), .ZN(n532) );
  XNOR2_X1 U626 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n533) );
  XOR2_X1 U627 ( .A(KEYINPUT100), .B(n534), .Z(n721) );
  NOR2_X1 U628 ( .A1(n721), .A2(n539), .ZN(n536) );
  XNOR2_X1 U629 ( .A(n536), .B(KEYINPUT31), .ZN(n698) );
  INV_X1 U630 ( .A(n580), .ZN(n537) );
  OR2_X1 U631 ( .A1(n537), .A2(n707), .ZN(n538) );
  NOR2_X1 U632 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U633 ( .A(KEYINPUT99), .B(n540), .Z(n541) );
  NAND2_X1 U634 ( .A1(n541), .A2(n579), .ZN(n686) );
  NAND2_X1 U635 ( .A1(n686), .A2(n698), .ZN(n546) );
  NOR2_X1 U636 ( .A1(n542), .A2(n545), .ZN(n543) );
  NAND2_X1 U637 ( .A1(n545), .A2(n542), .ZN(n696) );
  NAND2_X1 U638 ( .A1(n546), .A2(n596), .ZN(n547) );
  XNOR2_X1 U639 ( .A(n547), .B(KEYINPUT108), .ZN(n551) );
  NAND2_X1 U640 ( .A1(n605), .A2(n548), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n422), .A2(n549), .ZN(n550) );
  XNOR2_X1 U642 ( .A(n550), .B(KEYINPUT109), .ZN(n768) );
  INV_X1 U643 ( .A(n552), .ZN(n555) );
  INV_X1 U644 ( .A(n673), .ZN(n554) );
  NAND2_X1 U645 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U646 ( .A1(n556), .A2(KEYINPUT44), .ZN(n557) );
  XOR2_X1 U647 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n558) );
  NOR2_X1 U648 ( .A1(G900), .A2(n559), .ZN(n560) );
  NAND2_X1 U649 ( .A1(G953), .A2(n560), .ZN(n561) );
  XNOR2_X1 U650 ( .A(KEYINPUT111), .B(n561), .ZN(n564) );
  INV_X1 U651 ( .A(n562), .ZN(n563) );
  NOR2_X1 U652 ( .A1(n564), .A2(n563), .ZN(n600) );
  NAND2_X1 U653 ( .A1(n716), .A2(n399), .ZN(n567) );
  INV_X1 U654 ( .A(KEYINPUT30), .ZN(n566) );
  XNOR2_X1 U655 ( .A(n567), .B(n566), .ZN(n568) );
  BUF_X2 U656 ( .A(n570), .Z(n615) );
  INV_X1 U657 ( .A(KEYINPUT38), .ZN(n571) );
  XNOR2_X1 U658 ( .A(n615), .B(n571), .ZN(n724) );
  INV_X1 U659 ( .A(n724), .ZN(n572) );
  INV_X1 U660 ( .A(KEYINPUT39), .ZN(n573) );
  XNOR2_X1 U661 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n575) );
  XNOR2_X1 U662 ( .A(n576), .B(n575), .ZN(n766) );
  AND2_X1 U663 ( .A1(n713), .A2(n711), .ZN(n602) );
  INV_X1 U664 ( .A(n600), .ZN(n577) );
  NAND2_X1 U665 ( .A1(n602), .A2(n577), .ZN(n578) );
  XNOR2_X1 U666 ( .A(n580), .B(KEYINPUT113), .ZN(n581) );
  NOR2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n595) );
  INV_X1 U668 ( .A(n726), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n399), .A2(n583), .ZN(n584) );
  NOR2_X1 U670 ( .A1(n724), .A2(n584), .ZN(n586) );
  XNOR2_X1 U671 ( .A(KEYINPUT41), .B(KEYINPUT115), .ZN(n585) );
  NAND2_X1 U672 ( .A1(n595), .A2(n706), .ZN(n589) );
  XNOR2_X1 U673 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n587) );
  XNOR2_X1 U674 ( .A(n587), .B(KEYINPUT42), .ZN(n588) );
  XNOR2_X1 U675 ( .A(n589), .B(n588), .ZN(n767) );
  XNOR2_X1 U676 ( .A(n590), .B(KEYINPUT46), .ZN(n611) );
  NOR2_X1 U677 ( .A1(n591), .A2(n615), .ZN(n592) );
  XNOR2_X1 U678 ( .A(n592), .B(KEYINPUT112), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n594), .A2(n593), .ZN(n692) );
  NAND2_X1 U680 ( .A1(n595), .A2(n354), .ZN(n694) );
  XNOR2_X1 U681 ( .A(n597), .B(KEYINPUT47), .ZN(n598) );
  OR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U683 ( .A1(n696), .A2(n601), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n613) );
  NOR2_X1 U686 ( .A1(n613), .A2(n615), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n606), .B(KEYINPUT36), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n702) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT43), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n616), .A2(n394), .ZN(n704) );
  INV_X1 U692 ( .A(n704), .ZN(n617) );
  OR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  INV_X1 U694 ( .A(n620), .ZN(n703) );
  NAND2_X1 U695 ( .A1(n743), .A2(KEYINPUT2), .ZN(n621) );
  NOR2_X2 U696 ( .A1(n745), .A2(n621), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(n742) );
  NAND2_X1 U698 ( .A1(n743), .A2(n625), .ZN(n624) );
  OR2_X1 U699 ( .A1(n624), .A2(n745), .ZN(n629) );
  XOR2_X1 U700 ( .A(KEYINPUT81), .B(n625), .Z(n626) );
  NAND2_X1 U701 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  XOR2_X1 U702 ( .A(KEYINPUT69), .B(n627), .Z(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n742), .A2(n630), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n679), .A2(G472), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n637) );
  INV_X1 U707 ( .A(G952), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n635), .A2(G953), .ZN(n636) );
  NOR2_X2 U709 ( .A1(n637), .A2(n682), .ZN(n639) );
  INV_X1 U710 ( .A(KEYINPUT63), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(G57) );
  XNOR2_X1 U712 ( .A(n355), .B(G119), .ZN(G21) );
  XNOR2_X1 U713 ( .A(n641), .B(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n643), .B(n644), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT127), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n743), .B(n645), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n646), .A2(n473), .ZN(n651) );
  XNOR2_X1 U718 ( .A(n647), .B(G227), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n648), .A2(G900), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n649), .A2(G953), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(G72) );
  NAND2_X1 U722 ( .A1(n679), .A2(G475), .ZN(n655) );
  XNOR2_X1 U723 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U725 ( .A1(n656), .A2(n682), .ZN(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n679), .A2(G469), .ZN(n663) );
  BUF_X1 U729 ( .A(n659), .Z(n661) );
  XOR2_X1 U730 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n660) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X2 U732 ( .A1(n664), .A2(n682), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U734 ( .A1(n679), .A2(G210), .ZN(n670) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n667) );
  XNOR2_X1 U736 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X2 U737 ( .A1(n671), .A2(n682), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U739 ( .A(n673), .B(G122), .Z(G24) );
  BUF_X1 U740 ( .A(n679), .Z(n674) );
  NAND2_X1 U741 ( .A1(n674), .A2(G217), .ZN(n677) );
  BUF_X1 U742 ( .A(n675), .Z(n676) );
  XNOR2_X1 U743 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n678), .A2(n682), .ZN(G66) );
  NAND2_X1 U745 ( .A1(n674), .A2(G478), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(n680), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(G63) );
  NOR2_X1 U748 ( .A1(n686), .A2(n696), .ZN(n684) );
  XOR2_X1 U749 ( .A(G104), .B(n684), .Z(G6) );
  BUF_X1 U750 ( .A(n685), .Z(n699) );
  NOR2_X1 U751 ( .A1(n686), .A2(n699), .ZN(n688) );
  XNOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U754 ( .A(G107), .B(n689), .ZN(G9) );
  NOR2_X1 U755 ( .A1(n694), .A2(n699), .ZN(n691) );
  XNOR2_X1 U756 ( .A(G128), .B(KEYINPUT29), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n691), .B(n690), .ZN(G30) );
  XNOR2_X1 U758 ( .A(G143), .B(KEYINPUT118), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n693), .B(n692), .ZN(G45) );
  NOR2_X1 U760 ( .A1(n694), .A2(n696), .ZN(n695) );
  XOR2_X1 U761 ( .A(G146), .B(n695), .Z(G48) );
  NOR2_X1 U762 ( .A1(n696), .A2(n698), .ZN(n697) );
  XOR2_X1 U763 ( .A(G113), .B(n697), .Z(G15) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U765 ( .A(G116), .B(n700), .Z(G18) );
  XOR2_X1 U766 ( .A(G125), .B(KEYINPUT37), .Z(n701) );
  XNOR2_X1 U767 ( .A(n702), .B(n701), .ZN(G27) );
  XOR2_X1 U768 ( .A(G134), .B(n703), .Z(G36) );
  XNOR2_X1 U769 ( .A(n704), .B(G140), .ZN(n705) );
  XNOR2_X1 U770 ( .A(n705), .B(KEYINPUT119), .ZN(G42) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n710) );
  XOR2_X1 U772 ( .A(KEYINPUT121), .B(KEYINPUT50), .Z(n709) );
  XNOR2_X1 U773 ( .A(n710), .B(n709), .ZN(n719) );
  INV_X1 U774 ( .A(n711), .ZN(n712) );
  NAND2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U776 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n714) );
  XNOR2_X1 U777 ( .A(n715), .B(n714), .ZN(n717) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(KEYINPUT51), .B(n722), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n739), .A2(n723), .ZN(n734) );
  NOR2_X1 U783 ( .A1(n572), .A2(n399), .ZN(n725) );
  NOR2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U785 ( .A1(n572), .A2(n399), .ZN(n727) );
  NOR2_X1 U786 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n732) );
  INV_X1 U788 ( .A(n731), .ZN(n738) );
  NOR2_X1 U789 ( .A1(n732), .A2(n738), .ZN(n733) );
  NOR2_X1 U790 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U791 ( .A(n735), .B(KEYINPUT52), .ZN(n736) );
  NOR2_X1 U792 ( .A1(n737), .A2(n736), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n751) );
  NOR2_X1 U795 ( .A1(n743), .A2(KEYINPUT2), .ZN(n744) );
  XNOR2_X1 U796 ( .A(n744), .B(KEYINPUT80), .ZN(n748) );
  INV_X1 U797 ( .A(n745), .ZN(n754) );
  NOR2_X1 U798 ( .A1(n754), .A2(KEYINPUT2), .ZN(n746) );
  XOR2_X1 U799 ( .A(KEYINPUT79), .B(n746), .Z(n747) );
  NOR2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U801 ( .A1(n742), .A2(n749), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n752), .A2(G953), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n753), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U805 ( .A1(n754), .A2(n473), .ZN(n758) );
  NAND2_X1 U806 ( .A1(G953), .A2(G224), .ZN(n755) );
  XNOR2_X1 U807 ( .A(KEYINPUT61), .B(n755), .ZN(n756) );
  NAND2_X1 U808 ( .A1(n756), .A2(G898), .ZN(n757) );
  NAND2_X1 U809 ( .A1(n758), .A2(n757), .ZN(n765) );
  XOR2_X1 U810 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n763) );
  XOR2_X1 U811 ( .A(n759), .B(G101), .Z(n761) );
  OR2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n764) );
  XOR2_X1 U814 ( .A(n765), .B(n764), .Z(G69) );
  XOR2_X1 U815 ( .A(n766), .B(G131), .Z(G33) );
  XOR2_X1 U816 ( .A(n767), .B(G137), .Z(G39) );
  XNOR2_X1 U817 ( .A(G101), .B(n768), .ZN(G3) );
endmodule

