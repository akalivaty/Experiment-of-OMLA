//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1308,
    new_n1309, new_n1310, new_n1312, new_n1313, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0002(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n204));
  INV_X1    g0004(.A(G87), .ZN(new_n205));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n203), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  XOR2_X1   g0007(.A(KEYINPUT66), .B(G244), .Z(new_n208));
  AOI21_X1  g0008(.A(new_n207), .B1(G77), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  AOI22_X1  g0011(.A1(new_n209), .A2(new_n211), .B1(G1), .B2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT67), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n221), .B(new_n225), .C1(new_n212), .C2(new_n213), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n215), .A2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n218), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n219), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n247), .A2(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G50), .A2(G58), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n219), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n246), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT73), .B1(new_n219), .B2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT73), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G20), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G50), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n219), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n246), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n267), .B1(new_n263), .B2(new_n266), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT72), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(new_n246), .C1(new_n252), .C2(new_n255), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n257), .A2(new_n268), .A3(KEYINPUT9), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT74), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n257), .A2(new_n270), .A3(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n282), .A2(G223), .B1(new_n285), .B2(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n280), .A2(new_n281), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G1), .A3(G13), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n300), .A3(G274), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT70), .B1(new_n294), .B2(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G226), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n295), .A2(G190), .A3(new_n301), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n301), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n286), .B2(new_n292), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n276), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n273), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n312), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n271), .B(KEYINPUT74), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n295), .A2(new_n301), .A3(new_n307), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(G179), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n320), .A2(new_n274), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  XNOR2_X1  g0126(.A(G58), .B(G68), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n280), .A2(new_n219), .A3(new_n281), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n281), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT77), .B1(new_n333), .B2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n335), .B(new_n254), .C1(new_n331), .C2(new_n332), .ZN(new_n336));
  OAI211_X1 g0136(.A(KEYINPUT16), .B(new_n328), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT7), .B1(new_n285), .B2(new_n219), .ZN(new_n338));
  INV_X1    g0138(.A(new_n332), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n328), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n246), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n262), .A2(new_n247), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n267), .B1(new_n266), .B2(new_n247), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n300), .A2(G232), .A3(new_n304), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n301), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(G226), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G87), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n277), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n287), .C1(new_n283), .C2(new_n284), .ZN(new_n354));
  INV_X1    g0154(.A(G223), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n350), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n356), .B2(new_n294), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n321), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n359), .B(new_n349), .C1(new_n356), .C2(new_n294), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n326), .B1(new_n347), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n347), .A2(new_n326), .A3(new_n362), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(G190), .B2(new_n357), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(new_n344), .A3(new_n346), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n368), .A2(new_n344), .A3(KEYINPUT17), .A4(new_n346), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n364), .A2(new_n365), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n262), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(G77), .A3(new_n267), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n265), .A2(G1), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(G77), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G77), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n247), .A2(new_n251), .B1(new_n219), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n248), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n246), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n301), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n306), .B2(new_n208), .ZN(new_n387));
  INV_X1    g0187(.A(G232), .ZN(new_n388));
  INV_X1    g0188(.A(G107), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n354), .A2(new_n388), .B1(new_n389), .B2(new_n291), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(G238), .B2(new_n282), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(new_n300), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n392), .B2(new_n321), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n392), .A2(G179), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n385), .C1(new_n397), .C2(new_n392), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n325), .A2(new_n373), .A3(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n254), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n379), .B2(new_n248), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n246), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT11), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n266), .A2(new_n254), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT12), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(KEYINPUT11), .A3(new_n246), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n374), .A2(G68), .A3(new_n267), .ZN(new_n409));
  AND4_X1   g0209(.A1(new_n405), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n303), .B1(new_n300), .B2(new_n304), .ZN(new_n416));
  OAI21_X1  g0216(.A(G238), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n301), .ZN(new_n418));
  INV_X1    g0218(.A(G226), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n288), .A2(new_n289), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n388), .A2(new_n277), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n291), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n300), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n418), .A2(new_n424), .A3(KEYINPUT13), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n386), .B1(new_n306), .B2(G238), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n353), .A2(G226), .A3(new_n287), .ZN(new_n428));
  INV_X1    g0228(.A(new_n421), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n285), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n423), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n294), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n426), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n414), .B(G169), .C1(new_n425), .C2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT13), .B1(new_n418), .B2(new_n424), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n426), .A3(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(G179), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n414), .B1(new_n439), .B2(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n413), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n425), .A2(new_n433), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT14), .B1(new_n442), .B2(new_n321), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n437), .A4(new_n434), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n412), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(G200), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n412), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n400), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n219), .A2(G107), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n376), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT85), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT25), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n454), .A2(KEYINPUT25), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(KEYINPUT25), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n376), .A3(new_n452), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n246), .ZN(new_n459));
  OR3_X1    g0259(.A1(new_n279), .A2(KEYINPUT78), .A3(G1), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT78), .B1(new_n279), .B2(G1), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n459), .A2(new_n377), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n455), .B(new_n458), .C1(new_n462), .C2(new_n389), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G116), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n452), .A2(KEYINPUT23), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n219), .B2(G107), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n291), .A2(new_n219), .A3(G87), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(KEYINPUT22), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(KEYINPUT22), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT84), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n459), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n471), .B(KEYINPUT22), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n469), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT24), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n463), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G294), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n354), .C2(new_n206), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n290), .A2(G250), .A3(new_n291), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n485), .A4(new_n486), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n294), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n297), .A2(G1), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(G274), .A3(new_n300), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n300), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n502), .A2(G264), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n493), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT87), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n492), .B2(new_n294), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT87), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n496), .ZN(new_n509));
  AOI21_X1  g0309(.A(G190), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n366), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n484), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n480), .A2(KEYINPUT84), .A3(new_n477), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT24), .B1(new_n474), .B2(new_n475), .ZN(new_n515));
  AOI211_X1 g0315(.A(KEYINPUT84), .B(new_n470), .C1(new_n472), .C2(new_n473), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n246), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n463), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n508), .B1(new_n507), .B2(new_n496), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n300), .B1(new_n488), .B2(new_n491), .ZN(new_n521));
  INV_X1    g0321(.A(new_n496), .ZN(new_n522));
  NOR4_X1   g0322(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n522), .A4(new_n503), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n520), .A2(new_n523), .A3(new_n321), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n505), .A2(new_n359), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT82), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n250), .A2(G77), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n389), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  XNOR2_X1  g0332(.A(G97), .B(G107), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n529), .B1(new_n534), .B2(new_n219), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n389), .B1(new_n331), .B2(new_n332), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n246), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n266), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n462), .B2(new_n538), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G257), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n496), .B1(new_n501), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  INV_X1    g0345(.A(G244), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n354), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n282), .B2(G250), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT4), .A4(G244), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n544), .B1(new_n552), .B2(new_n294), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n321), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n359), .B(new_n544), .C1(new_n552), .C2(new_n294), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n542), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n548), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n354), .A2(new_n546), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(KEYINPUT4), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n300), .B1(new_n560), .B2(new_n547), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT80), .B(G200), .C1(new_n561), .C2(new_n544), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT80), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n553), .B2(new_n366), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  OAI21_X1  g0366(.A(G107), .B1(new_n338), .B2(new_n339), .ZN(new_n567));
  AND2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n532), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n530), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(G20), .B1(G77), .B2(new_n250), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n459), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n566), .B1(new_n573), .B2(new_n540), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n553), .A2(G190), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n537), .A2(KEYINPUT79), .A3(new_n541), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n556), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n579));
  INV_X1    g0379(.A(G238), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n464), .B(new_n579), .C1(new_n354), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n294), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n260), .A2(G45), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n300), .A2(G250), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n300), .A2(G274), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(new_n583), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n321), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n219), .B1(new_n423), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n569), .A2(new_n205), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n219), .B(G68), .C1(new_n283), .C2(new_n284), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n590), .B1(new_n248), .B2(new_n538), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n246), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n460), .A2(new_n461), .ZN(new_n598));
  INV_X1    g0398(.A(new_n381), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n267), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n381), .A2(new_n266), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n596), .A2(new_n246), .B1(new_n266), .B2(new_n381), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n586), .B1(new_n581), .B2(new_n294), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n359), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n589), .A2(new_n604), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n598), .A2(G87), .A3(new_n267), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(G190), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n612), .C1(new_n366), .C2(new_n607), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n528), .B1(new_n578), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n573), .A2(new_n566), .A3(new_n540), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT79), .B1(new_n537), .B2(new_n541), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n575), .A3(new_n564), .A4(new_n562), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n609), .A2(new_n613), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(KEYINPUT82), .A3(new_n556), .A4(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n548), .B(new_n219), .C1(G33), .C2(new_n538), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n622), .B(new_n246), .C1(new_n219), .C2(G116), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n266), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n598), .A2(G116), .A3(new_n267), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n500), .A2(G270), .A3(new_n300), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n496), .ZN(new_n631));
  OAI211_X1 g0431(.A(G264), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n280), .A2(G303), .A3(new_n281), .ZN(new_n633));
  OAI21_X1  g0433(.A(G257), .B1(new_n283), .B2(new_n284), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n353), .A2(new_n287), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n294), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n321), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT21), .B1(new_n629), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n637), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n397), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n366), .B1(new_n631), .B2(new_n637), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n629), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n630), .A2(new_n496), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n294), .B2(new_n636), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n638), .A2(KEYINPUT21), .B1(new_n646), .B2(G179), .ZN(new_n647));
  INV_X1    g0447(.A(new_n629), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(KEYINPUT21), .A3(G169), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(G179), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(KEYINPUT83), .A3(new_n629), .ZN(new_n653));
  AOI211_X1 g0453(.A(new_n639), .B(new_n643), .C1(new_n649), .C2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n615), .A2(new_n621), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n451), .A2(new_n527), .A3(new_n655), .ZN(G372));
  AND2_X1   g0456(.A1(new_n371), .A2(new_n372), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n412), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n321), .B1(new_n435), .B2(new_n436), .ZN(new_n660));
  AOI22_X1  g0460(.A1(G179), .A2(new_n442), .B1(new_n660), .B2(new_n414), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT76), .B1(new_n661), .B2(new_n443), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n438), .A2(new_n413), .A3(new_n440), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n448), .A2(new_n394), .A3(new_n393), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n658), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI211_X1 g0466(.A(KEYINPUT18), .B(new_n361), .C1(new_n344), .C2(new_n346), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n363), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT89), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n665), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n657), .B1(new_n445), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n668), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n318), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n588), .A2(new_n676), .A3(new_n321), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT88), .B1(new_n607), .B2(G169), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n602), .A4(new_n608), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n613), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  INV_X1    g0482(.A(new_n553), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G169), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n553), .A2(G179), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(new_n574), .B2(new_n576), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n542), .A3(new_n613), .A4(new_n609), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT26), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n690), .A3(new_n679), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n397), .B1(new_n520), .B2(new_n523), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n519), .B1(new_n692), .B2(new_n511), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n619), .A2(new_n681), .A3(new_n556), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n639), .B1(new_n629), .B2(new_n652), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n526), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n691), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n675), .B(new_n324), .C1(new_n451), .C2(new_n698), .ZN(G369));
  NAND2_X1  g0499(.A1(new_n376), .A2(new_n219), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT27), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G213), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(G343), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n513), .B(new_n526), .C1(new_n484), .C2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n506), .A2(G169), .A3(new_n509), .ZN(new_n709));
  INV_X1    g0509(.A(new_n525), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n484), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n706), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n706), .A2(new_n629), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT91), .ZN(new_n715));
  INV_X1    g0515(.A(new_n696), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n654), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n715), .ZN(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT92), .B(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n713), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n649), .A2(new_n653), .ZN(new_n724));
  INV_X1    g0524(.A(new_n639), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n706), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n513), .A2(new_n526), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n711), .A2(new_n707), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT93), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(KEYINPUT93), .A3(new_n728), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0534(.A(new_n223), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G41), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n592), .A2(G116), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n217), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n737), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n698), .B2(new_n706), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n578), .A2(new_n680), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n724), .A2(new_n725), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n513), .B(new_n745), .C1(new_n711), .C2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n679), .B1(new_n689), .B2(KEYINPUT26), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n682), .B1(new_n681), .B2(new_n686), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(KEYINPUT29), .A3(new_n707), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT96), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n744), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n615), .A2(new_n621), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n693), .A2(new_n711), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n756), .A3(new_n654), .A4(new_n707), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n640), .A2(new_n359), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n553), .A3(new_n607), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n493), .A2(new_n504), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n683), .A2(new_n588), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n763), .A2(KEYINPUT30), .A3(new_n507), .A4(new_n759), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n588), .A2(new_n640), .A3(new_n359), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT95), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n505), .A2(new_n683), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n762), .B(new_n764), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(KEYINPUT31), .B1(new_n769), .B2(new_n706), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n720), .B1(new_n757), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n706), .B1(new_n747), .B2(new_n750), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n754), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n742), .B1(new_n779), .B2(G1), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT97), .Z(G364));
  AND2_X1   g0581(.A1(new_n719), .A2(new_n721), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n265), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n260), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n736), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n721), .B2(new_n719), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n735), .A2(new_n285), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G355), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G116), .B2(new_n223), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n243), .A2(G45), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n735), .A2(new_n291), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n217), .B2(new_n297), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n218), .B1(G20), .B2(new_n321), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n786), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G179), .A2(G200), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n219), .B1(new_n804), .B2(G190), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT102), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT102), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G97), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n804), .A2(G20), .A3(new_n397), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G159), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n219), .A2(new_n366), .A3(G179), .A4(G190), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n816), .A2(KEYINPUT32), .B1(new_n818), .B2(new_n389), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n219), .A2(new_n359), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(G190), .A3(new_n366), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  INV_X1    g0622(.A(G58), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n820), .A2(new_n397), .A3(new_n366), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT99), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(KEYINPUT99), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n819), .B(new_n824), .C1(G77), .C2(new_n830), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n219), .A2(new_n397), .A3(new_n366), .A4(G179), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n285), .B1(new_n832), .B2(G87), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT100), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n820), .A2(G200), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n397), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(G190), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n263), .A2(new_n837), .B1(new_n839), .B2(new_n254), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(KEYINPUT32), .B2(new_n816), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n813), .A2(new_n831), .A3(new_n834), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G329), .ZN(new_n843));
  INV_X1    g0643(.A(G322), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n285), .B1(new_n814), .B2(new_n843), .C1(new_n821), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n830), .B2(G311), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n836), .A2(G326), .ZN(new_n847));
  XNOR2_X1  g0647(.A(KEYINPUT33), .B(G317), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n838), .A2(new_n848), .B1(G283), .B2(new_n817), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n832), .B(KEYINPUT103), .Z(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(G303), .ZN(new_n853));
  INV_X1    g0653(.A(G294), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n852), .A2(new_n853), .B1(new_n808), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n842), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n803), .B1(new_n856), .B2(new_n800), .ZN(new_n857));
  INV_X1    g0657(.A(new_n799), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n719), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n788), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G396));
  OAI211_X1 g0661(.A(new_n513), .B(new_n745), .C1(new_n711), .C2(new_n716), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n687), .A2(new_n690), .A3(new_n679), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n706), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n398), .B1(new_n385), .B2(new_n707), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n395), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n395), .A2(new_n706), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n864), .B(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n786), .B1(new_n871), .B2(new_n775), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n775), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n800), .A2(new_n797), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT104), .Z(new_n875));
  OAI21_X1  g0675(.A(new_n786), .B1(new_n875), .B2(G77), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT105), .Z(new_n877));
  INV_X1    g0677(.A(G283), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n878), .A2(new_n839), .B1(new_n837), .B2(new_n853), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G116), .B2(new_n830), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n818), .A2(new_n205), .ZN(new_n883));
  INV_X1    g0683(.A(G311), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n285), .B1(new_n814), .B2(new_n884), .C1(new_n821), .C2(new_n854), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n883), .B(new_n885), .C1(new_n851), .C2(G107), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n881), .A2(new_n813), .A3(new_n882), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n817), .A2(G68), .ZN(new_n888));
  INV_X1    g0688(.A(G132), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n888), .B(new_n291), .C1(new_n889), .C2(new_n814), .ZN(new_n890));
  INV_X1    g0690(.A(new_n808), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(G58), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n838), .A2(G150), .B1(new_n836), .B2(G137), .ZN(new_n893));
  INV_X1    g0693(.A(G143), .ZN(new_n894));
  INV_X1    g0694(.A(G159), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n893), .B1(new_n822), .B2(new_n894), .C1(new_n829), .C2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT34), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n892), .B1(new_n263), .B2(new_n852), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n887), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n877), .B1(new_n900), .B2(new_n800), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n870), .B2(new_n798), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n873), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(G384));
  OR2_X1    g0704(.A1(new_n571), .A2(KEYINPUT35), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n571), .A2(KEYINPUT35), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(G116), .A3(new_n220), .A4(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT36), .Z(new_n908));
  OAI211_X1 g0708(.A(new_n217), .B(G77), .C1(new_n823), .C2(new_n254), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n254), .A2(G50), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT107), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n260), .B(G13), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n757), .A2(new_n773), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n412), .A2(new_n707), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n664), .A2(new_n448), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT108), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n441), .A2(new_n444), .A3(new_n448), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n450), .A2(new_n918), .A3(new_n916), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n914), .A2(new_n870), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n347), .A2(new_n362), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n703), .A2(new_n705), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n347), .A2(new_n927), .ZN(new_n928));
  AND4_X1   g0728(.A1(new_n924), .A2(new_n925), .A3(new_n928), .A4(new_n369), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n337), .A2(new_n246), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n328), .B1(new_n334), .B2(new_n336), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT16), .B1(new_n931), .B2(KEYINPUT109), .ZN(new_n932));
  INV_X1    g0732(.A(new_n328), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n340), .A2(new_n335), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n333), .A2(KEYINPUT77), .A3(G68), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n930), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n346), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n927), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n362), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(new_n369), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n929), .B1(KEYINPUT37), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT38), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n657), .B2(new_n668), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n373), .A2(new_n347), .A3(new_n927), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n925), .A2(new_n928), .A3(new_n369), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT37), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n925), .A2(new_n928), .A3(new_n924), .A4(new_n369), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT38), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT40), .B1(new_n923), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n956));
  INV_X1    g0756(.A(new_n941), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n373), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n369), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n459), .B1(new_n936), .B2(KEYINPUT16), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n342), .B1(new_n936), .B2(new_n937), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n931), .A2(KEYINPUT109), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n346), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n959), .B1(new_n964), .B2(new_n362), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n924), .B1(new_n965), .B2(new_n941), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n958), .B(KEYINPUT38), .C1(new_n966), .C2(new_n929), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT40), .B1(new_n956), .B2(new_n967), .ZN(new_n968));
  NOR4_X1   g0768(.A1(new_n445), .A2(KEYINPUT108), .A3(new_n449), .A4(new_n915), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n917), .B2(new_n920), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n869), .B1(new_n757), .B2(new_n773), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n955), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n914), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n451), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n720), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n956), .A2(KEYINPUT39), .A3(new_n967), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n950), .A2(new_n951), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n928), .B1(new_n657), .B2(new_n668), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n945), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT39), .B1(new_n981), .B2(new_n967), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n445), .A2(new_n707), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n864), .A2(new_n870), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n868), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n956), .A2(new_n967), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n989), .A3(new_n970), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n669), .A2(new_n926), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n451), .B1(new_n754), .B2(new_n777), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n675), .A2(new_n324), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n992), .B(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n977), .A2(new_n996), .B1(new_n260), .B2(new_n783), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n977), .A2(new_n996), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n913), .B1(new_n997), .B2(new_n998), .ZN(G367));
  OAI221_X1 g0799(.A(new_n801), .B1(new_n223), .B2(new_n381), .C1(new_n234), .C2(new_n794), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(new_n786), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n707), .A2(new_n611), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n681), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n679), .B2(new_n1002), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n839), .A2(new_n895), .B1(new_n379), .B2(new_n818), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n291), .B1(new_n249), .B2(new_n821), .C1(new_n837), .C2(new_n894), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G50), .C2(new_n830), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n812), .A2(G68), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n832), .A2(G58), .B1(new_n815), .B2(G137), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT113), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n285), .B1(new_n814), .B2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n854), .A2(new_n839), .B1(new_n837), .B2(new_n884), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G97), .C2(new_n817), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n851), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n389), .C2(new_n808), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT46), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n832), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n626), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n822), .B2(new_n853), .C1(new_n829), .C2(new_n878), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1011), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  INV_X1    g0823(.A(new_n800), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1001), .B1(new_n858), .B2(new_n1004), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n726), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n708), .A2(new_n712), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n727), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n782), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n722), .A2(new_n1027), .A3(new_n727), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1031), .A2(new_n754), .A3(new_n775), .A4(new_n777), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n619), .B(new_n556), .C1(new_n618), .C2(new_n707), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n686), .A2(new_n706), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n727), .A2(KEYINPUT93), .A3(new_n728), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT93), .B1(new_n727), .B2(new_n728), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT45), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(KEYINPUT45), .B(new_n1035), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1035), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n731), .A2(new_n1043), .A3(new_n732), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT44), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n731), .A2(new_n1043), .A3(KEYINPUT44), .A4(new_n732), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n723), .A2(KEYINPUT111), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1032), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1041), .A2(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n1050), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n778), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n736), .B(KEYINPUT41), .Z(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT112), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n778), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1053), .B2(new_n1050), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n779), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1056), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n785), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1043), .A2(new_n727), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT42), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(KEYINPUT42), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n556), .B1(new_n1043), .B2(new_n526), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1068), .A2(new_n1069), .B1(new_n707), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1071), .A2(KEYINPUT110), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT110), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(new_n1072), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1073), .A2(new_n1074), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n723), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n1043), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1077), .B(new_n1079), .Z(new_n1080));
  OAI21_X1  g0880(.A(new_n1025), .B1(new_n1066), .B2(new_n1080), .ZN(G387));
  NAND2_X1  g0881(.A1(new_n778), .A2(new_n1058), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n1032), .A3(new_n736), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n713), .A2(new_n799), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n738), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(new_n789), .B1(new_n389), .B2(new_n735), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n231), .A2(new_n297), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n247), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n263), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT50), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n738), .B(new_n297), .C1(new_n254), .C2(new_n379), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n793), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n801), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n811), .A2(new_n381), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n836), .A2(G159), .B1(G97), .B2(new_n817), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n838), .A2(new_n1088), .B1(G77), .B2(new_n832), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n291), .B1(new_n814), .B2(new_n249), .C1(new_n821), .C2(new_n263), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n830), .B2(G68), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT114), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n808), .A2(new_n878), .B1(new_n854), .B2(new_n1019), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n838), .A2(G311), .B1(new_n836), .B2(G322), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n822), .B2(new_n1012), .C1(new_n829), .C2(new_n853), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT48), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT49), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n291), .B1(new_n815), .B2(G326), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n626), .B2(new_n818), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1109), .B2(KEYINPUT49), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1102), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n786), .B(new_n1094), .C1(new_n1114), .C2(new_n1024), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1083), .B1(new_n784), .B2(new_n1058), .C1(new_n1084), .C2(new_n1115), .ZN(G393));
  AOI21_X1  g0916(.A(new_n737), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1053), .B(new_n1078), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT116), .B1(new_n1118), .B2(new_n1032), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1049), .A2(new_n723), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1053), .A2(new_n1078), .ZN(new_n1121));
  OAI211_X1 g0921(.A(KEYINPUT116), .B(new_n1032), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1117), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1118), .A2(new_n784), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1043), .A2(new_n799), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n239), .A2(new_n793), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n801), .B1(new_n538), .B2(new_n223), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n786), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n285), .B1(new_n814), .B2(new_n844), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n839), .A2(new_n853), .B1(new_n878), .B2(new_n1019), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(G107), .C2(new_n817), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n837), .A2(new_n1012), .B1(new_n884), .B2(new_n821), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n891), .A2(G116), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n830), .A2(G294), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n837), .A2(new_n249), .B1(new_n895), .B2(new_n821), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT51), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n839), .A2(new_n263), .B1(new_n254), .B2(new_n1019), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n291), .B1(new_n814), .B2(new_n894), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1140), .A2(new_n883), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(new_n247), .C2(new_n829), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n811), .A2(new_n379), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1129), .B1(new_n1145), .B2(new_n800), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1125), .B1(new_n1126), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1124), .A2(new_n1147), .ZN(G390));
  NOR3_X1   g0948(.A1(new_n655), .A2(new_n527), .A3(new_n706), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n772), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n770), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n870), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n921), .A2(new_n922), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n706), .B(new_n869), .C1(new_n862), .C2(new_n863), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n921), .B(new_n922), .C1(new_n1155), .C2(new_n867), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT39), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n947), .B2(new_n953), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n956), .A2(new_n967), .A3(KEYINPUT39), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1156), .A2(new_n984), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n867), .B1(new_n776), .B2(new_n866), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(new_n1153), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n981), .A2(new_n967), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n984), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1154), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n984), .B(new_n1163), .C1(new_n1161), .C2(new_n1153), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n970), .A2(new_n774), .A3(new_n870), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n985), .B1(new_n988), .B2(new_n970), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1168), .C1(new_n983), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n774), .A2(new_n870), .B1(new_n921), .B2(new_n922), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n988), .B1(new_n1172), .B2(new_n1154), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1168), .A2(new_n1161), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(G330), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n974), .A2(new_n1177), .A3(new_n451), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n993), .A2(new_n994), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n737), .B1(new_n1171), .B2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1166), .A2(new_n1176), .A3(new_n1170), .A4(new_n1179), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n786), .B1(new_n875), .B2(new_n1088), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n291), .B1(new_n851), .B2(G87), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n888), .B1(new_n626), .B2(new_n821), .C1(new_n854), .C2(new_n814), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n389), .A2(new_n839), .B1(new_n837), .B2(new_n878), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(G97), .C2(new_n830), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(new_n1189), .C1(new_n379), .C2(new_n811), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT119), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n830), .A2(new_n1193), .B1(G137), .B2(new_n838), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n811), .B2(new_n895), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT117), .Z(new_n1196));
  NAND2_X1  g0996(.A1(new_n832), .A2(G150), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT53), .Z(new_n1198));
  NOR2_X1   g0998(.A1(new_n821), .A2(new_n889), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n285), .B(new_n1199), .C1(G125), .C2(new_n815), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n836), .A2(G128), .B1(G50), .B2(new_n817), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1191), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1184), .B1(new_n1203), .B2(new_n800), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n983), .B2(new_n798), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1171), .B2(new_n784), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1183), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(G378));
  AND3_X1   g1008(.A1(new_n986), .A2(new_n990), .A3(new_n991), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT122), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n927), .A2(new_n1210), .A3(new_n274), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n927), .B2(new_n274), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n325), .A2(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1215));
  INV_X1    g1015(.A(new_n1213), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n318), .A2(new_n324), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1215), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n323), .B(new_n1213), .C1(new_n313), .C2(new_n317), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n318), .B2(new_n324), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n973), .B2(G330), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1218), .A2(new_n1222), .A3(KEYINPUT123), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT123), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1177), .B(new_n1228), .C1(new_n955), .C2(new_n972), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1209), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n970), .A2(new_n1163), .A3(new_n971), .ZN(new_n1231));
  AND4_X1   g1031(.A1(new_n914), .A2(new_n870), .A3(new_n921), .A4(new_n922), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1231), .A2(KEYINPUT40), .B1(new_n1232), .B2(new_n968), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1223), .B1(new_n1233), .B2(new_n1177), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1228), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n973), .A2(G330), .A3(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n992), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n784), .B1(new_n1230), .B2(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n538), .A2(new_n839), .B1(new_n837), .B2(new_n626), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1019), .A2(new_n379), .B1(new_n818), .B2(new_n823), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n291), .A2(G41), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n878), .B2(new_n814), .C1(new_n389), .C2(new_n821), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n830), .B2(new_n599), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1008), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT58), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G50), .B(new_n1242), .C1(new_n279), .C2(new_n296), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT120), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT121), .B1(new_n832), .B2(new_n1193), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n832), .A2(KEYINPUT121), .A3(new_n1193), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n830), .C2(G137), .ZN(new_n1253));
  INV_X1    g1053(.A(G128), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n839), .A2(new_n889), .B1(new_n1254), .B2(new_n821), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G125), .B2(new_n836), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1253), .B(new_n1256), .C1(new_n249), .C2(new_n811), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n817), .A2(G159), .ZN(new_n1260));
  AOI211_X1 g1060(.A(G33), .B(G41), .C1(new_n815), .C2(G124), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1250), .B1(KEYINPUT58), .B2(new_n1246), .C1(new_n1258), .C2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n800), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n786), .C1(G50), .C2(new_n875), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1235), .B2(new_n797), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1238), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1182), .A2(new_n1179), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1182), .A2(KEYINPUT124), .A3(new_n1179), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT57), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1230), .B2(new_n1237), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1182), .A2(KEYINPUT124), .A3(new_n1179), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT124), .B1(new_n1182), .B2(new_n1179), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n736), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1267), .B1(new_n1274), .B2(new_n1280), .ZN(G375));
  OR3_X1    g1081(.A1(new_n993), .A2(new_n994), .A3(new_n1178), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1064), .A3(new_n1180), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1176), .A2(new_n785), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n970), .A2(new_n798), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n291), .B1(new_n814), .B2(new_n1254), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n889), .A2(new_n837), .B1(new_n839), .B2(new_n1192), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(G58), .C2(new_n817), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n822), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n830), .A2(G150), .B1(new_n1290), .B2(G137), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1289), .B(new_n1291), .C1(new_n895), .C2(new_n852), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n811), .A2(new_n263), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n839), .A2(new_n626), .B1(new_n379), .B2(new_n818), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(G294), .B2(new_n836), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n851), .A2(G97), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n830), .A2(G107), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n285), .B1(new_n821), .B2(new_n878), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(G303), .B2(new_n815), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .A4(new_n1299), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n1292), .A2(new_n1293), .B1(new_n1300), .B2(new_n1095), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n800), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1302), .B(new_n786), .C1(G68), .C2(new_n875), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1286), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1285), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1284), .A2(new_n1306), .ZN(G381));
  AND2_X1   g1107(.A1(new_n1124), .A2(new_n1147), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1308), .A2(new_n1306), .A3(new_n1284), .A4(new_n1309), .ZN(new_n1310));
  OR4_X1    g1110(.A1(G387), .A2(G375), .A3(new_n1310), .A4(G378), .ZN(G407));
  NOR2_X1   g1111(.A1(new_n704), .A2(G343), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1207), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G407), .B(G213), .C1(G375), .C2(new_n1313), .ZN(G409));
  NAND2_X1  g1114(.A1(G387), .A2(new_n1308), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G390), .B(new_n1025), .C1(new_n1066), .C2(new_n1080), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(G393), .B(new_n860), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT127), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1180), .A2(new_n736), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT125), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1283), .A2(new_n1327), .A3(KEYINPUT60), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT60), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1326), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(G384), .A3(new_n1306), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n903), .B1(new_n1332), .B2(new_n1305), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1312), .A2(G2897), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1336), .B(new_n1337), .ZN(new_n1338));
  OAI211_X1 g1138(.A(G378), .B(new_n1267), .C1(new_n1274), .C2(new_n1280), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1267), .B1(new_n1340), .B2(new_n1056), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1207), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1312), .B1(new_n1339), .B2(new_n1342), .ZN(new_n1343));
  AOI211_X1 g1143(.A(new_n1312), .B(new_n1336), .C1(new_n1339), .C2(new_n1342), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  OAI221_X1 g1145(.A(new_n1325), .B1(new_n1338), .B2(new_n1343), .C1(new_n1344), .C2(new_n1345), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1324), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1312), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1335), .ZN(new_n1350));
  OR2_X1    g1150(.A1(new_n1238), .A2(new_n1266), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n737), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1340), .A2(new_n1275), .ZN(new_n1353));
  AOI211_X1 g1153(.A(new_n1207), .B(new_n1351), .C1(new_n1352), .C2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1342), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1349), .B(new_n1350), .C1(new_n1354), .C2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1320), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1336), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT63), .B1(new_n1343), .B2(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1325), .B1(new_n1338), .B2(new_n1343), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT126), .B1(new_n1360), .B2(new_n1362), .ZN(new_n1363));
  OAI211_X1 g1163(.A(new_n1356), .B(new_n1320), .C1(new_n1344), .C2(KEYINPUT63), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT126), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1364), .A2(new_n1365), .A3(new_n1361), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1348), .B1(new_n1363), .B2(new_n1366), .ZN(G405));
  AND2_X1   g1167(.A1(G375), .A2(new_n1207), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1368), .A2(new_n1354), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1336), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1358), .B1(new_n1368), .B2(new_n1354), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  XNOR2_X1  g1172(.A(new_n1372), .B(new_n1324), .ZN(G402));
endmodule


