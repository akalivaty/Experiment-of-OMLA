//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n205), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n215), .B1(new_n216), .B2(new_n205), .C1(new_n217), .C2(new_n212), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR4_X1   g0026(.A1(new_n218), .A2(new_n220), .A3(new_n223), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT64), .B(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G238), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n208), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT1), .Z(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n202), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n214), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n225), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  INV_X1    g0049(.A(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(KEYINPUT66), .B(G107), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n248), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G232), .A3(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT72), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n266), .A3(G232), .A4(G1698), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n261), .A2(new_n264), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n255), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n268), .A2(new_n271), .B1(G238), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI211_X1 g0082(.A(G1), .B(new_n277), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n275), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n276), .B1(new_n275), .B2(new_n284), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT14), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n286), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n275), .A2(new_n276), .A3(new_n284), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(G169), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n289), .B(new_n294), .C1(new_n295), .C2(new_n292), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT73), .B(KEYINPUT12), .Z(new_n297));
  NAND2_X1  g0097(.A1(new_n206), .A2(G20), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT69), .B1(new_n298), .B2(new_n209), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n207), .A2(G1), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(G13), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n297), .B1(new_n303), .B2(new_n228), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT74), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n303), .A2(KEYINPUT12), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(G68), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n299), .A2(new_n302), .ZN(new_n308));
  NAND3_X1  g0108(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n232), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n308), .A2(new_n310), .A3(new_n300), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT68), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n309), .A2(new_n314), .A3(new_n232), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G20), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G50), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n207), .A2(G33), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n319), .B1(new_n221), .B2(new_n320), .C1(new_n228), .C2(new_n207), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT11), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n307), .A2(new_n312), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n296), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n260), .A2(G232), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT70), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n262), .A2(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G238), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n217), .B2(new_n262), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n271), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n274), .A2(G244), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n284), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n288), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n311), .A2(G77), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT15), .B(G87), .Z(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n320), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT8), .B(G58), .ZN(new_n339));
  INV_X1    g0139(.A(new_n318), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(new_n207), .B2(new_n221), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n310), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n335), .B(new_n342), .C1(G77), .C2(new_n303), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n334), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n333), .A2(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n324), .B1(new_n292), .B2(G200), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n287), .A2(G190), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n325), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n317), .A2(new_n308), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(G50), .A3(new_n298), .ZN(new_n352));
  INV_X1    g0152(.A(G50), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n207), .B1(new_n201), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G150), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n339), .A2(new_n320), .B1(new_n355), .B2(new_n340), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n317), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n352), .B(new_n357), .C1(G50), .C2(new_n303), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT9), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n259), .A2(new_n221), .ZN(new_n360));
  MUX2_X1   g0160(.A(G222), .B(G223), .S(G1698), .Z(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n271), .C1(new_n259), .C2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G226), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n284), .B(new_n362), .C1(new_n363), .C2(new_n273), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G200), .B2(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n368), .B(new_n371), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n364), .A2(G179), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n364), .A2(new_n288), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n358), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n339), .A2(new_n300), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n351), .A2(new_n377), .B1(new_n308), .B2(new_n339), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n310), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n257), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT7), .B(new_n207), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n262), .B2(G20), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n259), .A2(KEYINPUT77), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n228), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n340), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n201), .B1(new_n228), .B2(G58), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n391), .B(new_n394), .C1(new_n395), .C2(new_n207), .ZN(new_n396));
  INV_X1    g0196(.A(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT64), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT64), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G68), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n400), .A3(G58), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n207), .B1(new_n401), .B2(new_n202), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT75), .B1(new_n402), .B2(new_n393), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n390), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n380), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n387), .A2(new_n383), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n403), .A2(new_n396), .A3(KEYINPUT76), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT76), .B1(new_n403), .B2(new_n396), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT16), .B(new_n408), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n379), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n363), .A2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n262), .B(new_n413), .C1(G223), .C2(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n283), .B1(new_n416), .B2(new_n271), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n274), .A2(G232), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G200), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G190), .B2(new_n419), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n412), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n422), .ZN(new_n426));
  INV_X1    g0226(.A(new_n390), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n403), .A2(new_n396), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n405), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n411), .A2(new_n310), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n378), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n419), .A2(new_n295), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n288), .B1(new_n417), .B2(new_n418), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT18), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n412), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n425), .B(new_n426), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n343), .B1(new_n333), .B2(G200), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n365), .B2(new_n333), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n350), .A2(new_n376), .A3(new_n439), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n308), .A2(new_n219), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n206), .A2(G33), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n351), .A2(G97), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n389), .A2(KEYINPUT79), .A3(G107), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT79), .B1(new_n389), .B2(G107), .ZN(new_n449));
  XNOR2_X1  g0249(.A(G97), .B(G107), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT6), .A2(G107), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G20), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n221), .B2(new_n340), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n448), .A2(new_n449), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n444), .B(new_n446), .C1(new_n458), .C2(new_n380), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n206), .B(G45), .C1(new_n460), .C2(G41), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT67), .B(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n463), .A2(new_n211), .A3(new_n271), .ZN(new_n464));
  INV_X1    g0264(.A(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n262), .A2(G244), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT4), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n465), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n464), .B1(new_n472), .B2(new_n271), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n463), .A2(G274), .ZN(new_n474));
  AOI21_X1  g0274(.A(G169), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(new_n277), .A3(new_n461), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n464), .B(new_n477), .C1(new_n472), .C2(new_n271), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n295), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n459), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n389), .A2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT79), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n447), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n310), .B1(new_n484), .B2(new_n457), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n473), .A2(new_n365), .A3(new_n474), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n478), .B2(G200), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n485), .A2(new_n487), .A3(new_n444), .A4(new_n446), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n262), .A2(new_n207), .A3(G68), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n320), .B2(new_n219), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n207), .B1(new_n265), .B2(new_n490), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT80), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n207), .C1(new_n265), .C2(new_n490), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NOR4_X1   g0296(.A1(KEYINPUT81), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT81), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n216), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n489), .B(new_n491), .C1(new_n496), .C2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n310), .B1(new_n308), .B2(new_n337), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n351), .A2(new_n336), .A3(new_n445), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n329), .A2(new_n465), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n222), .A2(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n256), .A2(new_n505), .A3(new_n258), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n270), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n206), .A2(G45), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n270), .A2(G250), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n277), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n503), .A2(new_n504), .B1(new_n515), .B2(new_n288), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n295), .ZN(new_n517));
  NOR4_X1   g0317(.A1(new_n509), .A2(new_n512), .A3(new_n365), .A4(new_n513), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n515), .B2(G200), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n502), .A2(new_n310), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n308), .A2(new_n337), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n316), .A2(new_n303), .A3(G87), .A4(new_n445), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n516), .A2(new_n517), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n480), .A2(new_n488), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT82), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT82), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n480), .A2(new_n488), .A3(new_n527), .A4(new_n524), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n256), .A2(new_n258), .A3(G257), .A4(new_n465), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n256), .A2(new_n258), .A3(G264), .A4(G1698), .ZN(new_n530));
  INV_X1    g0330(.A(G303), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n262), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n271), .ZN(new_n533));
  OAI211_X1 g0333(.A(G270), .B(new_n270), .C1(new_n476), .C2(new_n461), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n474), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n250), .B1(new_n206), .B2(G33), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n303), .A2(new_n380), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n299), .A2(new_n302), .A3(new_n250), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n250), .A2(G20), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n310), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n471), .B(new_n207), .C1(G33), .C2(new_n219), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT20), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND4_X1   g0343(.A1(KEYINPUT20), .A2(new_n542), .A3(new_n310), .A4(new_n540), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n538), .B(new_n539), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n536), .B(new_n546), .C1(new_n365), .C2(new_n535), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT83), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n535), .A2(new_n545), .A3(G169), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n535), .A2(new_n295), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n535), .A2(new_n545), .A3(KEYINPUT21), .A4(G169), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n260), .A2(G250), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n211), .C2(new_n328), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n271), .ZN(new_n560));
  OAI211_X1 g0360(.A(G264), .B(new_n270), .C1(new_n476), .C2(new_n461), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n560), .A2(new_n474), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n295), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT25), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n308), .A2(new_n564), .A3(new_n217), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n316), .A2(new_n303), .A3(G107), .A4(new_n445), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT25), .B1(new_n303), .B2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT85), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT85), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n262), .A2(new_n207), .A3(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n262), .A2(new_n575), .A3(new_n207), .A4(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(KEYINPUT23), .A2(G107), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(G20), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(KEYINPUT84), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(KEYINPUT84), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n577), .A2(KEYINPUT24), .A3(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n310), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n572), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n560), .A2(new_n474), .A3(new_n561), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n288), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n563), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n562), .A2(G190), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(G200), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n572), .A3(new_n589), .A4(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n548), .A2(new_n556), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n443), .A2(new_n526), .A3(new_n528), .A4(new_n597), .ZN(G372));
  NAND2_X1  g0398(.A1(new_n516), .A2(new_n517), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n459), .A2(new_n479), .A3(new_n524), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT26), .ZN(new_n602));
  XNOR2_X1  g0402(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n459), .A2(new_n524), .A3(new_n479), .A4(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n480), .A2(new_n488), .A3(new_n524), .A4(new_n596), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n555), .A2(KEYINPUT86), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT86), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n551), .A2(new_n553), .A3(new_n608), .A4(new_n554), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n607), .A2(new_n593), .A3(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n602), .B(new_n605), .C1(new_n606), .C2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n443), .B1(new_n600), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n375), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n325), .A2(new_n346), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n422), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT17), .B1(new_n412), .B2(new_n422), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n617), .A3(new_n349), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n431), .A2(new_n435), .A3(KEYINPUT18), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n437), .B1(new_n412), .B2(new_n434), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n613), .B1(new_n622), .B2(new_n372), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n612), .A2(new_n623), .ZN(G369));
  NOR2_X1   g0424(.A1(new_n209), .A2(G20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n206), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT89), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n548), .B(new_n556), .C1(new_n546), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n607), .A2(new_n609), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n545), .A3(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n590), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n596), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n593), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n593), .A2(new_n633), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n556), .A2(new_n633), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT90), .B1(new_n648), .B2(new_n643), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(KEYINPUT90), .A3(new_n643), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n649), .B2(new_n651), .ZN(G399));
  NAND2_X1  g0452(.A1(new_n501), .A2(new_n250), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n210), .A2(new_n462), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(G1), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n234), .B2(new_n656), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT28), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n601), .A2(new_n604), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n459), .A2(new_n524), .A3(KEYINPUT26), .A4(new_n479), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n600), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n663), .B2(new_n662), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n593), .A2(new_n556), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n606), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n663), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n600), .B1(new_n670), .B2(KEYINPUT92), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT93), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n667), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(KEYINPUT29), .A3(new_n634), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n634), .B1(new_n611), .B2(new_n600), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT91), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT91), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n679), .B(new_n634), .C1(new_n611), .C2(new_n600), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n526), .A2(new_n597), .A3(new_n528), .A4(new_n634), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n562), .A2(new_n473), .A3(new_n514), .A4(new_n552), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT30), .Z(new_n685));
  INV_X1    g0485(.A(new_n478), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n535), .ZN(new_n687));
  NOR4_X1   g0487(.A1(new_n687), .A2(G179), .A3(new_n514), .A4(new_n562), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n633), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n689), .A2(KEYINPUT31), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n682), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n659), .B1(new_n695), .B2(G1), .ZN(G364));
  INV_X1    g0496(.A(new_n638), .ZN(new_n697));
  NOR2_X1   g0497(.A1(G13), .A2(G33), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G20), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n625), .A2(G45), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n656), .A2(G1), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n210), .A2(new_n262), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n248), .B2(G45), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G45), .B2(new_n234), .ZN(new_n708));
  INV_X1    g0508(.A(new_n210), .ZN(new_n709));
  INV_X1    g0509(.A(G355), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n262), .ZN(new_n711));
  OAI221_X1 g0511(.A(new_n708), .B1(G116), .B2(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n232), .B1(G20), .B2(new_n288), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n700), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n207), .A2(G190), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n420), .A2(G179), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n217), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G159), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n207), .A2(new_n365), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n717), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n723), .A2(KEYINPUT32), .B1(new_n216), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n295), .A2(new_n420), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n719), .B(new_n726), .C1(G50), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n295), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n716), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G77), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n723), .A2(KEYINPUT32), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n724), .A2(new_n731), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n207), .B1(new_n720), .B2(G190), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n224), .B1(new_n737), .B2(new_n219), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n727), .A2(new_n716), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n259), .B(new_n738), .C1(G68), .C2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n730), .A2(new_n734), .A3(new_n735), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G326), .ZN(new_n743));
  INV_X1    g0543(.A(G311), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n728), .A2(new_n743), .B1(new_n732), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n737), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(G294), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  INV_X1    g0548(.A(new_n718), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G283), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n262), .B1(new_n722), .B2(G329), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  INV_X1    g0552(.A(new_n725), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n740), .A2(new_n752), .B1(new_n753), .B2(G303), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G322), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n736), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n742), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n713), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n701), .A2(new_n704), .A3(new_n715), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n697), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n639), .A3(new_n703), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(G396));
  NOR2_X1   g0564(.A1(new_n346), .A2(new_n633), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n633), .A2(new_n343), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n441), .A2(new_n766), .B1(new_n344), .B2(new_n345), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n677), .A2(new_n680), .A3(new_n769), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n768), .B(new_n634), .C1(new_n600), .C2(new_n611), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(new_n693), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n693), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n773), .A2(new_n703), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n698), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n753), .B1(new_n749), .B2(G68), .ZN(new_n777));
  INV_X1    g0577(.A(new_n736), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G143), .A2(new_n778), .B1(new_n733), .B2(G159), .ZN(new_n779));
  INV_X1    g0579(.A(G137), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n779), .B1(new_n780), .B2(new_n728), .C1(new_n355), .C2(new_n739), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n262), .B(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  INV_X1    g0584(.A(G132), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n785), .B2(new_n721), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n783), .B(new_n786), .C1(G58), .C2(new_n746), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G116), .A2(new_n733), .B1(new_n722), .B2(G311), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n788), .B1(new_n217), .B2(new_n725), .C1(new_n531), .C2(new_n728), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n259), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n718), .A2(new_n216), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n736), .A2(new_n796), .B1(new_n737), .B2(new_n219), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n789), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n713), .B1(new_n787), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n713), .A2(new_n698), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n221), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n776), .A2(new_n704), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n775), .A2(new_n802), .ZN(G384));
  AND3_X1   g0603(.A1(new_n296), .A2(new_n324), .A3(new_n634), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n324), .A2(new_n633), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n296), .A2(new_n324), .B1(new_n349), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND4_X1   g0607(.A1(new_n690), .A2(new_n807), .A3(new_n691), .A4(new_n768), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n411), .A2(new_n317), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n405), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n379), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n423), .B1(new_n812), .B2(new_n631), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n434), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT37), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n431), .B1(new_n435), .B2(new_n630), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT37), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n816), .A2(new_n817), .A3(new_n423), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT97), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n811), .A2(new_n411), .A3(new_n317), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n378), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n630), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(new_n617), .C2(new_n621), .ZN(new_n824));
  INV_X1    g0624(.A(new_n823), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT97), .B1(new_n439), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(KEYINPUT38), .B(new_n819), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n816), .A2(new_n423), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(new_n817), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n412), .B(new_n631), .C1(new_n617), .C2(new_n621), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n808), .A2(new_n833), .A3(KEYINPUT40), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT98), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n439), .A2(new_n825), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n820), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n439), .A2(KEYINPUT97), .A3(new_n825), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n839), .B2(new_n819), .ZN(new_n840));
  INV_X1    g0640(.A(new_n827), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n819), .B1(new_n824), .B2(new_n826), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n828), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(KEYINPUT98), .A3(new_n827), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(new_n845), .A3(new_n808), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT40), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n834), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n443), .A3(new_n692), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n761), .B(new_n834), .C1(new_n846), .C2(new_n847), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n692), .A2(new_n443), .A3(G330), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n675), .A2(new_n681), .A3(new_n443), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n623), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n853), .B(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n765), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n771), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n807), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n842), .A2(new_n860), .A3(new_n845), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n833), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n844), .A2(KEYINPUT39), .A3(new_n827), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n804), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n619), .A2(new_n620), .A3(new_n631), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n861), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n856), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n206), .B2(new_n625), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n250), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n871), .B(new_n233), .C1(KEYINPUT35), .C2(new_n455), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n235), .A2(G77), .A3(new_n401), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(G50), .B2(new_n397), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(G1), .A3(new_n209), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n873), .A3(new_n876), .ZN(G367));
  AOI22_X1  g0677(.A1(G283), .A2(new_n733), .B1(new_n722), .B2(G317), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n749), .A2(G97), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n878), .B(new_n879), .C1(new_n744), .C2(new_n728), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(G303), .B2(new_n778), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n725), .A2(new_n250), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n882), .A2(KEYINPUT46), .B1(new_n217), .B2(new_n737), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n262), .B(new_n883), .C1(KEYINPUT46), .C2(new_n882), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n881), .B(new_n884), .C1(new_n796), .C2(new_n792), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT106), .Z(new_n886));
  OAI21_X1  g0686(.A(new_n262), .B1(new_n792), .B2(new_n392), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G68), .B2(new_n746), .ZN(new_n888));
  AOI22_X1  g0688(.A1(G50), .A2(new_n733), .B1(new_n749), .B2(G77), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n780), .B2(new_n721), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G143), .B2(new_n729), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n753), .A2(G58), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n778), .A2(G150), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n888), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT47), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n713), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n714), .B1(new_n709), .B2(new_n337), .C1(new_n243), .C2(new_n706), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n704), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n634), .A2(new_n523), .ZN(new_n900));
  MUX2_X1   g0700(.A(new_n524), .B(new_n600), .S(new_n900), .Z(new_n901));
  NOR3_X1   g0701(.A1(new_n901), .A2(G20), .A3(new_n699), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n655), .B(KEYINPUT41), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n639), .A2(KEYINPUT105), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n639), .B2(KEYINPUT105), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n648), .A2(KEYINPUT104), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n695), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n649), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n459), .A2(new_n633), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n480), .A2(new_n915), .A3(new_n488), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n459), .A2(new_n479), .A3(new_n633), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(new_n650), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n914), .A2(KEYINPUT44), .A3(new_n650), .A4(new_n919), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(KEYINPUT102), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n918), .B1(new_n651), .B2(new_n649), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT45), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(KEYINPUT45), .B(new_n918), .C1(new_n651), .C2(new_n649), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT102), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n920), .A2(new_n930), .A3(new_n921), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n645), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n924), .A2(new_n929), .A3(new_n646), .A4(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n905), .B(new_n913), .C1(new_n935), .C2(KEYINPUT103), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n904), .B1(new_n936), .B2(new_n694), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n702), .A2(G1), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n919), .A2(new_n648), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(KEYINPUT101), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(KEYINPUT101), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n918), .B(KEYINPUT100), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n480), .B1(new_n946), .B2(new_n593), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n634), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n944), .B1(new_n942), .B2(new_n943), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n901), .B(KEYINPUT99), .Z(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n950), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n646), .A2(new_n946), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n903), .B1(new_n940), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(G387));
  AOI22_X1  g0761(.A1(G317), .A2(new_n778), .B1(new_n733), .B2(G303), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n756), .B2(new_n728), .C1(new_n792), .C2(new_n744), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT48), .Z(new_n964));
  OAI22_X1  g0764(.A1(new_n725), .A2(new_n796), .B1(new_n737), .B2(new_n793), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT110), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT110), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n259), .B1(new_n968), .B2(KEYINPUT49), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT49), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n250), .B2(new_n718), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(G326), .C2(new_n722), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n337), .A2(new_n737), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n732), .A2(new_n397), .B1(new_n721), .B2(new_n355), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n778), .A2(G50), .ZN(new_n976));
  INV_X1    g0776(.A(new_n339), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n740), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n975), .A2(new_n879), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n725), .A2(new_n221), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n728), .A2(new_n392), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n979), .A2(new_n259), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n713), .B1(new_n972), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n644), .A2(new_n700), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n240), .A2(new_n282), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n653), .A2(KEYINPUT108), .ZN(new_n990));
  AOI21_X1  g0790(.A(G45), .B1(new_n653), .B2(KEYINPUT108), .ZN(new_n991));
  NAND2_X1  g0791(.A1(G68), .A2(G77), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n339), .A2(G50), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n988), .A2(new_n989), .A3(new_n705), .A4(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(G107), .B2(new_n709), .C1(new_n654), .C2(new_n711), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n703), .B(new_n985), .C1(new_n714), .C2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n912), .B2(new_n938), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n913), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n655), .B1(new_n695), .B2(new_n912), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(G393));
  NAND2_X1  g0803(.A1(new_n935), .A2(new_n913), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n1001), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n655), .B(new_n1004), .C1(new_n1006), .C2(new_n905), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n933), .A2(new_n938), .A3(new_n934), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n946), .A2(new_n700), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G317), .A2(new_n729), .B1(new_n778), .B2(G311), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT52), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n259), .B1(new_n793), .B2(new_n725), .C1(new_n792), .C2(new_n531), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n719), .B(new_n1012), .C1(G322), .C2(new_n722), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n746), .A2(G116), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1011), .B(new_n1015), .C1(G294), .C2(new_n733), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n753), .A2(new_n228), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n262), .B(new_n1017), .C1(new_n792), .C2(new_n353), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n977), .B2(new_n733), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n746), .A2(G77), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n728), .A2(new_n355), .B1(new_n736), .B2(new_n392), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT51), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n795), .B1(G143), .B2(new_n722), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT111), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n713), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n253), .A2(new_n705), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n714), .C1(new_n219), .C2(new_n709), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1009), .A2(new_n704), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1007), .A2(new_n1008), .A3(new_n1029), .ZN(G390));
  NAND4_X1  g0830(.A1(new_n690), .A2(new_n807), .A3(new_n691), .A4(new_n768), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n761), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n804), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n833), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n806), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n767), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n674), .A2(new_n634), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n857), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1034), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n863), .A2(new_n864), .B1(new_n1033), .B2(new_n859), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n863), .A2(new_n864), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n859), .A2(new_n1033), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1038), .A2(new_n1035), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1034), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n808), .A2(G330), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n854), .A2(new_n623), .A3(new_n851), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n690), .A2(new_n691), .A3(G330), .A4(new_n768), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n807), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n858), .B1(new_n1054), .B2(new_n1032), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1048), .A2(new_n857), .A3(new_n1037), .A4(new_n1053), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1041), .A2(new_n1049), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n655), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1041), .A2(new_n1049), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1057), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1042), .A2(new_n698), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n718), .A2(new_n397), .B1(new_n721), .B2(new_n796), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT113), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n792), .A2(new_n217), .B1(new_n793), .B2(new_n728), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n778), .A2(G116), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n262), .B1(new_n746), .B2(G77), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G87), .A2(new_n753), .B1(new_n733), .B2(G97), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT54), .B(G143), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n732), .A2(new_n1072), .B1(new_n737), .B2(new_n392), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n792), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(G137), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT112), .Z(new_n1076));
  AOI22_X1  g0876(.A1(G50), .A2(new_n749), .B1(new_n722), .B2(G125), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n753), .A2(G150), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT53), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n259), .B(new_n1079), .C1(G128), .C2(new_n729), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n736), .A2(new_n785), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1071), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n713), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n800), .A2(new_n339), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1063), .A2(new_n704), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1060), .B2(new_n939), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1062), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G378));
  INV_X1    g0889(.A(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n358), .A2(new_n630), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n376), .B(new_n1091), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n850), .B2(KEYINPUT117), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n867), .B1(new_n850), .B2(KEYINPUT117), .ZN(new_n1099));
  AND4_X1   g0899(.A1(KEYINPUT117), .A2(new_n848), .A3(G330), .A4(new_n867), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n848), .A2(G330), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT117), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1096), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n850), .A2(KEYINPUT117), .A3(new_n867), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n848), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n868), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1050), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1058), .A2(KEYINPUT118), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT118), .B1(new_n1058), .B2(new_n1110), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1090), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1058), .A2(new_n1110), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1058), .A2(KEYINPUT118), .A3(new_n1110), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(KEYINPUT57), .A3(new_n1108), .A4(new_n1101), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1114), .A2(new_n655), .A3(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n713), .A2(G50), .A3(new_n698), .ZN(new_n1122));
  INV_X1    g0922(.A(G124), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n255), .B(new_n269), .C1(new_n721), .C2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n739), .A2(new_n785), .B1(new_n732), .B2(new_n780), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G128), .B2(new_n778), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n729), .A2(G125), .B1(new_n746), .B2(G150), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n725), .C2(new_n1072), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT59), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1124), .B(new_n1129), .C1(G159), .C2(new_n749), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n262), .A2(new_n462), .ZN(new_n1131));
  AOI211_X1 g0931(.A(G50), .B(new_n1131), .C1(new_n255), .C2(new_n269), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1131), .B1(new_n221), .B2(new_n725), .C1(new_n219), .C2(new_n739), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n778), .A2(G107), .B1(new_n746), .B2(G68), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n722), .A2(G283), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n749), .A2(G58), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n733), .A2(new_n336), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1133), .B(new_n1138), .C1(G116), .C2(new_n729), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n1140));
  XNOR2_X1  g0940(.A(new_n1139), .B(new_n1140), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1130), .A2(new_n1132), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n703), .B(new_n1122), .C1(new_n1143), .C2(new_n713), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1097), .B2(new_n699), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1109), .B2(new_n939), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1121), .A2(new_n1147), .ZN(G375));
  AOI21_X1  g0948(.A(new_n939), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1052), .A2(new_n698), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n725), .A2(new_n219), .B1(new_n721), .B2(new_n531), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT119), .Z(new_n1152));
  AOI22_X1  g0952(.A1(G107), .A2(new_n733), .B1(new_n749), .B2(G77), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n259), .C1(new_n793), .C2(new_n736), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n792), .A2(new_n250), .B1(new_n796), .B2(new_n728), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .A4(new_n973), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n792), .A2(new_n1072), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n259), .B1(new_n746), .B2(G50), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n753), .A2(G159), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n778), .A2(G137), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1136), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n722), .A2(G128), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n728), .A2(new_n785), .B1(new_n732), .B2(new_n355), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1157), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n713), .B1(new_n1156), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n800), .A2(new_n397), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1150), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1149), .B1(new_n704), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1055), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n904), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1170), .B2(new_n1057), .ZN(G381));
  NOR2_X1   g0971(.A1(G375), .A2(G378), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(G390), .A2(G381), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G387), .B1(KEYINPUT120), .B2(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(KEYINPUT120), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .A4(new_n1177), .ZN(G407));
  NAND2_X1  g0978(.A1(new_n632), .A2(G213), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1172), .A2(KEYINPUT121), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(G407), .A2(G213), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT121), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1182), .A2(new_n1183), .ZN(G409));
  INV_X1    g0984(.A(KEYINPUT61), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1121), .A2(G378), .A3(new_n1147), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n904), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1109), .A2(new_n1113), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1088), .B1(new_n1188), .B2(new_n1146), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1180), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n656), .B1(new_n1169), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1061), .C1(new_n1191), .C2(new_n1169), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1193), .A2(G384), .A3(new_n1168), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G384), .B1(new_n1193), .B2(new_n1168), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1180), .A2(G2897), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1185), .B1(new_n1190), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT124), .ZN(new_n1200));
  INV_X1    g1000(.A(G390), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(G387), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(G393), .B(G396), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT122), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n960), .B2(G390), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n940), .A2(new_n959), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n903), .ZN(new_n1207));
  INV_X1    g1007(.A(G396), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(G393), .B(new_n1208), .ZN(new_n1209));
  AND4_X1   g1009(.A1(new_n1206), .A2(new_n1207), .A3(G390), .A4(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1202), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(G387), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n1185), .C1(new_n1190), .C2(new_n1198), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1200), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT62), .Z(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT63), .B1(new_n1190), .B2(new_n1198), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1217), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1221), .A2(KEYINPUT63), .A3(new_n1179), .A4(new_n1196), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT123), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT123), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1190), .A2(new_n1224), .A3(KEYINPUT63), .A4(new_n1196), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1185), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1216), .A2(new_n1218), .B1(new_n1226), .B2(new_n1227), .ZN(G405));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(KEYINPUT126), .B(KEYINPUT127), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1213), .A2(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1186), .A2(KEYINPUT125), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1196), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1186), .A2(KEYINPUT125), .A3(new_n1196), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n1088), .A3(G375), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G375), .A2(new_n1088), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1238), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1196), .B1(new_n1186), .B2(KEYINPUT125), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1233), .A2(new_n1234), .A3(new_n1239), .A4(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1234), .A2(new_n1243), .A3(new_n1239), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(G402));
endmodule


