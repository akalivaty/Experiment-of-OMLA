//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n208), .A2(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  AND3_X1   g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT64), .B(G238), .Z(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT65), .Z(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n216), .B1(new_n209), .B2(new_n208), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT67), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G1), .ZN(new_n247));
  AND3_X1   g0047(.A1(new_n245), .A2(new_n247), .A3(G20), .ZN(new_n248));
  OR2_X1    g0048(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT67), .B(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n213), .B1(new_n206), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n249), .A2(new_n250), .A3(new_n252), .A4(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n260), .A2(KEYINPUT73), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(KEYINPUT73), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT15), .B(G87), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n214), .A2(G33), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(new_n214), .B2(new_n257), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n254), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G77), .B2(new_n252), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n213), .ZN(new_n270));
  AND3_X1   g0070(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT66), .B1(G33), .B2(G41), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n245), .B(new_n247), .C1(G41), .C2(G45), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G244), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI211_X1 g0079(.A(G1), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT72), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G107), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n286), .A2(new_n222), .B1(new_n287), .B2(new_n285), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G232), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n292), .A2(new_n293), .A3(G1698), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n284), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(G200), .B1(new_n283), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n276), .B2(new_n281), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n297), .B(new_n295), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n269), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n283), .B2(new_n295), .ZN(new_n305));
  OAI211_X1 g0105(.A(G179), .B(new_n295), .C1(new_n298), .C2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n303), .B1(new_n308), .B2(new_n269), .ZN(new_n309));
  INV_X1    g0109(.A(new_n252), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(G50), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n256), .B2(G50), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT8), .A2(G58), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT69), .B(G58), .Z(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(KEYINPUT8), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(new_n214), .A3(G33), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n255), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n285), .A2(G222), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n323), .B1(new_n257), .B2(new_n285), .C1(new_n286), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n284), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n280), .B1(new_n275), .B2(G226), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n321), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n321), .A3(new_n327), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n320), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n330), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n332), .A2(new_n328), .A3(new_n304), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n319), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT71), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(KEYINPUT71), .B(new_n319), .C1(new_n331), .C2(new_n333), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n309), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  OR2_X1    g0139(.A1(KEYINPUT79), .A2(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(KEYINPUT79), .A2(G33), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT3), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n291), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT7), .B(new_n214), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n285), .B2(G20), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n221), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n201), .B1(new_n314), .B2(G68), .ZN(new_n348));
  INV_X1    g0148(.A(G159), .ZN(new_n349));
  INV_X1    g0149(.A(new_n260), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n348), .A2(new_n214), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n339), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT69), .B(G58), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n210), .B1(new_n353), .B2(new_n221), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n340), .A2(KEYINPUT3), .A3(new_n341), .ZN(new_n356));
  AOI21_X1  g0156(.A(G20), .B1(new_n356), .B2(new_n290), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n357), .B2(new_n345), .ZN(new_n358));
  AOI211_X1 g0158(.A(KEYINPUT7), .B(G20), .C1(new_n356), .C2(new_n290), .ZN(new_n359));
  OAI211_X1 g0159(.A(KEYINPUT16), .B(new_n355), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n352), .A2(new_n360), .A3(new_n254), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n273), .A2(new_n274), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n281), .B1(new_n363), .B2(new_n293), .ZN(new_n364));
  INV_X1    g0164(.A(new_n284), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G226), .A2(G1698), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n324), .B2(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n290), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n362), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n275), .A2(G232), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n368), .A2(new_n369), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(new_n281), .C1(new_n373), .C2(new_n365), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n371), .B1(new_n374), .B2(G190), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n256), .A2(new_n315), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n310), .B2(new_n315), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n361), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n361), .A2(new_n377), .A3(new_n375), .A4(KEYINPUT17), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n304), .B1(new_n364), .B2(new_n370), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n374), .B2(G179), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n361), .B2(new_n377), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI211_X1 g0187(.A(KEYINPUT18), .B(new_n384), .C1(new_n361), .C2(new_n377), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n382), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT74), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n312), .A2(new_n318), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(KEYINPUT9), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT9), .ZN(new_n393));
  NOR4_X1   g0193(.A1(new_n312), .A2(new_n318), .A3(KEYINPUT74), .A4(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n319), .A2(new_n393), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n329), .A2(G200), .A3(new_n330), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT10), .ZN(new_n399));
  OAI21_X1  g0199(.A(G190), .B1(new_n332), .B2(new_n328), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n395), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n400), .A3(new_n397), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n392), .A2(new_n394), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT10), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n338), .A2(new_n389), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n310), .A2(new_n254), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(G68), .A3(new_n249), .A4(new_n250), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n257), .B2(new_n265), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n410), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT11), .B1(new_n410), .B2(new_n254), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OR3_X1    g0213(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n408), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT76), .B(KEYINPUT13), .Z(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n290), .A2(new_n291), .A3(G226), .A4(new_n322), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n290), .A2(new_n291), .A3(G232), .A4(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(KEYINPUT75), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n284), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n273), .A2(new_n274), .A3(G238), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n281), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n419), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n427), .A3(new_n419), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n304), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n426), .A2(new_n281), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n285), .A2(new_n438), .A3(G232), .A4(G1698), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n437), .A2(new_n439), .A3(new_n420), .A4(new_n421), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n284), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n430), .B(G179), .C1(new_n435), .C2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n431), .B2(new_n432), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n418), .B1(new_n434), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n430), .B(G190), .C1(new_n435), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n417), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n425), .A2(new_n427), .A3(new_n419), .ZN(new_n447));
  OAI21_X1  g0247(.A(G200), .B1(new_n447), .B2(new_n428), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT77), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(G200), .C1(new_n447), .C2(new_n428), .ZN(new_n451));
  AOI211_X1 g0251(.A(KEYINPUT78), .B(new_n446), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT78), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n451), .ZN(new_n454));
  INV_X1    g0254(.A(new_n446), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n444), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n406), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n340), .A2(new_n341), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n343), .B1(new_n459), .B2(new_n289), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n346), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G107), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n350), .A2(new_n257), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT6), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n465), .A2(new_n466), .B1(new_n469), .B2(G107), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n287), .A2(G97), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n473));
  OAI211_X1 g0273(.A(G97), .B(new_n287), .C1(new_n467), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n464), .B1(new_n475), .B2(G20), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI211_X1 g0278(.A(KEYINPUT81), .B(new_n464), .C1(new_n475), .C2(G20), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n254), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n251), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n252), .A2(new_n481), .A3(G97), .A4(new_n255), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G97), .B2(new_n252), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT82), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n245), .A2(new_n247), .A3(G45), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(new_n273), .A3(G274), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n251), .A2(new_n488), .A3(G45), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n273), .ZN(new_n491));
  INV_X1    g0291(.A(G257), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n322), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n356), .A2(G244), .A3(new_n322), .A4(new_n290), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n499), .A2(KEYINPUT83), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT83), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n493), .B1(new_n503), .B2(new_n284), .ZN(new_n504));
  OR3_X1    g0304(.A1(new_n504), .A2(KEYINPUT84), .A3(new_n362), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT84), .B1(new_n504), .B2(new_n362), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n486), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(G190), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT85), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n504), .A2(new_n304), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n320), .B(new_n493), .C1(new_n503), .C2(new_n284), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n486), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n264), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n252), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n214), .B1(new_n516), .B2(new_n420), .ZN(new_n517));
  INV_X1    g0317(.A(G87), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n469), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(G107), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n221), .A2(G20), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n356), .A2(new_n290), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT87), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT87), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n356), .A2(new_n524), .A3(new_n290), .A4(new_n521), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n516), .B1(G20), .B2(new_n420), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n520), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n515), .B1(new_n527), .B2(new_n254), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n407), .A2(new_n481), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n514), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n356), .A2(G238), .A3(new_n322), .A4(new_n290), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n356), .A2(G244), .A3(G1698), .A4(new_n290), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n459), .A2(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n245), .A2(new_n247), .A3(G45), .A4(new_n277), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n273), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n487), .A2(G250), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n535), .A2(new_n284), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G179), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n304), .B2(new_n540), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n297), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G200), .B2(new_n540), .ZN(new_n544));
  AND4_X1   g0344(.A1(G87), .A2(new_n252), .A3(new_n255), .A4(new_n481), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n515), .B(new_n545), .C1(new_n527), .C2(new_n254), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n531), .A2(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n513), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(G264), .A2(G1698), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n356), .A2(new_n290), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT88), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n292), .A2(G303), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n356), .A2(G257), .A3(new_n322), .A4(new_n290), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n356), .A2(KEYINPUT88), .A3(new_n290), .A4(new_n550), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n284), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n490), .A2(G270), .A3(new_n273), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n489), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n252), .A2(new_n481), .A3(G116), .A4(new_n255), .ZN(new_n563));
  INV_X1    g0363(.A(G116), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n248), .A2(G13), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n253), .A2(G97), .ZN(new_n567));
  AOI21_X1  g0367(.A(G20), .B1(new_n567), .B2(new_n496), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n214), .A2(new_n564), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n254), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(KEYINPUT20), .B(new_n254), .C1(new_n568), .C2(new_n569), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n304), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n562), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n566), .A2(new_n574), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n562), .A2(G190), .ZN(new_n581));
  AOI21_X1  g0381(.A(G200), .B1(new_n558), .B2(new_n561), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n562), .A2(KEYINPUT21), .A3(new_n575), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT89), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n579), .A2(new_n558), .A3(G179), .A4(new_n561), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n578), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n287), .A3(G20), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT90), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n214), .A2(G87), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n292), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n356), .A2(KEYINPUT22), .A3(G87), .A4(new_n290), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n534), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n214), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(G20), .B1(new_n600), .B2(new_n534), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT24), .B1(new_n605), .B2(new_n598), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT91), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(new_n602), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT91), .B1(new_n609), .B2(KEYINPUT24), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n254), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n529), .A2(G107), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT25), .B1(new_n252), .B2(G107), .ZN(new_n613));
  OR3_X1    g0413(.A1(new_n252), .A2(KEYINPUT25), .A3(G107), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n490), .A2(G264), .A3(new_n273), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n322), .A2(G250), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n492), .B2(new_n322), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n356), .A2(new_n620), .A3(new_n290), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n459), .A2(G294), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n365), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n489), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n297), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G200), .B2(new_n625), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n611), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n609), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n606), .A2(new_n607), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n604), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n615), .B1(new_n631), .B2(new_n254), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n625), .A2(new_n304), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(G179), .B2(new_n625), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n628), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n589), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n458), .A2(new_n510), .A3(new_n549), .A4(new_n636), .ZN(G372));
  XNOR2_X1  g0437(.A(new_n385), .B(KEYINPUT18), .ZN(new_n638));
  INV_X1    g0438(.A(new_n444), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n452), .A2(new_n456), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n308), .A2(new_n269), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n638), .B1(new_n642), .B2(new_n382), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n405), .B1(new_n336), .B2(new_n337), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n584), .A2(new_n586), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n645), .B(new_n578), .C1(new_n632), .C2(new_n634), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n510), .A2(new_n549), .A3(new_n628), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n542), .A2(new_n531), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n544), .A2(new_n546), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n513), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n493), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n499), .A2(new_n500), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT83), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n499), .A2(KEYINPUT83), .A3(new_n500), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n497), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n658), .B2(new_n365), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G169), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n504), .A2(G179), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n660), .A2(new_n661), .B1(new_n485), .B2(new_n480), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n547), .A3(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n652), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n647), .A2(new_n648), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n458), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n644), .A2(new_n666), .ZN(G369));
  AND2_X1   g0467(.A1(new_n214), .A2(G13), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n251), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n628), .B1(new_n632), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n632), .A2(new_n634), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n632), .A2(new_n634), .A3(new_n674), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT93), .Z(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n580), .A2(new_n675), .ZN(new_n683));
  INV_X1    g0483(.A(new_n589), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n685), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n645), .A2(new_n578), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n683), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n682), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n587), .ZN(new_n692));
  INV_X1    g0492(.A(new_n588), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n577), .B2(new_n576), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n674), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n681), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n696), .A3(new_n679), .ZN(G399));
  INV_X1    g0497(.A(new_n207), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n519), .A2(G107), .A3(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n211), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n548), .B1(new_n507), .B2(new_n509), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n636), .A2(new_n705), .A3(new_n675), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n320), .B(new_n560), .C1(new_n557), .C2(new_n284), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n504), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT94), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n618), .A2(new_n623), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n540), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n709), .B1(new_n540), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n708), .A2(KEYINPUT30), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n540), .A2(new_n710), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT94), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n540), .A2(new_n710), .A3(new_n709), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n504), .A3(new_n707), .A4(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n625), .A2(new_n540), .A3(G179), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n659), .A3(new_n562), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n674), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n722), .B1(new_n718), .B2(new_n719), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT30), .B1(new_n708), .B2(new_n713), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT31), .B(new_n674), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n706), .B1(new_n730), .B2(KEYINPUT95), .ZN(new_n731));
  INV_X1    g0531(.A(new_n729), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n723), .B2(new_n674), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT95), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n665), .A2(new_n675), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n663), .A2(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n663), .A2(KEYINPUT96), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT97), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n652), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT97), .B(new_n649), .C1(new_n513), .C2(new_n651), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n743), .A2(new_n744), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n694), .A2(new_n677), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n705), .A3(new_n628), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n750), .A3(new_n648), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n739), .B1(new_n742), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n704), .B1(new_n753), .B2(G1), .ZN(G364));
  NAND3_X1  g0554(.A1(new_n687), .A2(new_n682), .A3(new_n689), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n690), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(KEYINPUT98), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n668), .A2(G45), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n700), .A2(G1), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n756), .B2(KEYINPUT98), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n687), .A2(new_n689), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n213), .B1(G20), .B2(new_n304), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n214), .A2(new_n297), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n320), .A2(new_n362), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n292), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n214), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(G329), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n320), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n774), .B(new_n779), .C1(G322), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n776), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G294), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n362), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n770), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT100), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G303), .ZN(new_n791));
  XOR2_X1   g0591(.A(KEYINPUT33), .B(G317), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n771), .A2(new_n775), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n775), .A2(new_n787), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n775), .A2(new_n780), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G311), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n783), .A2(new_n786), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n772), .A2(new_n202), .B1(new_n781), .B2(new_n353), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n292), .B(new_n801), .C1(G77), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n785), .A2(G97), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n777), .A2(new_n349), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n794), .A2(new_n287), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n788), .A2(new_n518), .ZN(new_n808));
  INV_X1    g0608(.A(new_n793), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n808), .C1(G68), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n802), .A2(new_n803), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n769), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n766), .A2(new_n768), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n356), .A2(new_n290), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n698), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n239), .A2(new_n279), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n212), .A2(G45), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n698), .A2(new_n292), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G355), .B1(new_n564), .B2(new_n698), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n761), .B(new_n812), .C1(new_n813), .C2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n759), .A2(new_n763), .B1(new_n767), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n768), .A2(new_n764), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n761), .B1(new_n257), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n794), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G87), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n292), .ZN(new_n830));
  INV_X1    g0630(.A(new_n772), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G303), .B1(new_n778), .B2(G311), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n564), .B2(new_n797), .C1(new_n795), .C2(new_n793), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n830), .B(new_n833), .C1(G107), .C2(new_n790), .ZN(new_n834));
  INV_X1    g0634(.A(G294), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n803), .B1(new_n835), .B2(new_n781), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT101), .Z(new_n837));
  AOI22_X1  g0637(.A1(new_n831), .A2(G137), .B1(new_n798), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G143), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n839), .B2(new_n781), .C1(new_n840), .C2(new_n793), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT34), .ZN(new_n842));
  INV_X1    g0642(.A(new_n785), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n353), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n815), .B1(new_n221), .B2(new_n794), .C1(new_n845), .C2(new_n777), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(G50), .C2(new_n790), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n834), .A2(new_n837), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n641), .A2(new_n675), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n674), .B1(new_n258), .B2(new_n268), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n303), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n851), .B2(new_n641), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n827), .B1(new_n769), .B2(new_n848), .C1(new_n853), .C2(new_n765), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n740), .B(new_n853), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n762), .B1(new_n739), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n739), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(G384));
  INV_X1    g0659(.A(KEYINPUT104), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n361), .A2(new_n377), .ZN(new_n862));
  INV_X1    g0662(.A(new_n384), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n672), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n866), .A3(new_n378), .ZN(new_n867));
  XNOR2_X1  g0667(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n864), .A2(new_n866), .A3(new_n378), .A4(new_n868), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n380), .A2(new_n381), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n866), .B1(new_n638), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n860), .B(new_n861), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n339), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n254), .A3(new_n360), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(new_n377), .B1(new_n384), .B2(new_n672), .ZN(new_n879));
  INV_X1    g0679(.A(new_n378), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n871), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n377), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n865), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT38), .B(new_n882), .C1(new_n389), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n870), .A2(new_n871), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n389), .B2(new_n866), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n860), .B1(new_n888), .B2(new_n861), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n417), .A2(new_n675), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n457), .A2(new_n891), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n444), .B1(new_n417), .B2(new_n675), .C1(new_n452), .C2(new_n456), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n852), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n734), .A2(new_n706), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT40), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n884), .B1(new_n638), .B2(new_n873), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n881), .A2(new_n871), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n861), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n885), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(new_n901), .A3(new_n895), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT106), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n897), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n458), .A2(new_n895), .ZN(new_n910));
  OAI21_X1  g0710(.A(G330), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n752), .A2(new_n458), .A3(new_n742), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n752), .A2(new_n742), .A3(KEYINPUT105), .A4(new_n458), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n915), .A2(new_n644), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n901), .A2(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n638), .A2(new_n873), .ZN(new_n919));
  INV_X1    g0719(.A(new_n866), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n919), .A2(new_n920), .B1(new_n871), .B2(new_n870), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT104), .B1(new_n921), .B2(KEYINPUT38), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n885), .A3(new_n875), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n923), .B2(KEYINPUT39), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n444), .A2(new_n674), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n638), .A2(new_n865), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n892), .A2(new_n893), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n665), .A2(new_n853), .A3(new_n675), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n849), .B(KEYINPUT102), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n927), .B1(new_n932), .B2(new_n901), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n917), .B(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n912), .A2(new_n935), .B1(new_n251), .B2(new_n668), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n912), .B2(new_n935), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n212), .B(G77), .C1(new_n221), .C2(new_n353), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n202), .A2(G68), .ZN(new_n939));
  AOI211_X1 g0739(.A(G13), .B(new_n251), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(G116), .B(new_n215), .C1(new_n475), .C2(KEYINPUT35), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(KEYINPUT35), .B2(new_n475), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n937), .A2(new_n940), .A3(new_n943), .ZN(G367));
  AOI21_X1  g0744(.A(new_n662), .B1(new_n486), .B2(new_n674), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n510), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n662), .A2(new_n674), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n946), .A2(new_n677), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n674), .B1(new_n951), .B2(new_n513), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT42), .B1(new_n696), .B2(new_n949), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n546), .A2(new_n675), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n547), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n648), .A2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n953), .A2(new_n954), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n691), .A2(new_n949), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n691), .B2(new_n949), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n699), .B(KEYINPUT41), .Z(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n696), .A2(new_n679), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n968), .B1(new_n970), .B2(new_n948), .ZN(new_n971));
  INV_X1    g0771(.A(new_n968), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n949), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n969), .B2(new_n949), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n696), .A2(KEYINPUT45), .A3(new_n679), .A4(new_n948), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n691), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n973), .A3(new_n971), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n690), .A3(new_n681), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n681), .B(new_n695), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n690), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n753), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n979), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n967), .B1(new_n986), .B2(new_n753), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n760), .A2(G1), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n964), .B(new_n966), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n816), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n813), .B1(new_n207), .B2(new_n264), .C1(new_n990), .C2(new_n235), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n762), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n790), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G283), .A2(new_n798), .B1(new_n778), .B2(G317), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G294), .A2(new_n809), .B1(new_n782), .B2(G303), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n788), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT46), .B1(new_n997), .B2(G116), .ZN(new_n998));
  INV_X1    g0798(.A(G311), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n814), .B1(new_n469), .B2(new_n794), .C1(new_n999), .C2(new_n772), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(G107), .C2(new_n785), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n772), .A2(new_n839), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n793), .A2(new_n349), .B1(new_n797), .B2(new_n202), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(G150), .C2(new_n782), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n828), .A2(G77), .ZN(new_n1005));
  INV_X1    g0805(.A(G137), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n777), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n843), .A2(new_n221), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n788), .A2(new_n353), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n292), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n996), .A2(new_n1001), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n769), .B1(new_n1011), .B2(KEYINPUT47), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n992), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n766), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n958), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n989), .A2(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n983), .A2(new_n988), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n997), .A2(G294), .B1(new_n785), .B2(G283), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n831), .A2(G322), .B1(new_n798), .B2(G303), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n999), .B2(new_n793), .C1(new_n1021), .C2(new_n781), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT49), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n794), .A2(new_n564), .B1(new_n777), .B2(new_n773), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1026), .A2(new_n815), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G159), .A2(new_n831), .B1(new_n997), .B2(G77), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n782), .B1(new_n798), .B2(G68), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n315), .A2(new_n809), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n843), .A2(new_n264), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n794), .A2(new_n469), .B1(new_n777), .B2(new_n840), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1032), .A2(new_n814), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n768), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n259), .A2(G50), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT50), .Z(new_n1038));
  OAI211_X1 g0838(.A(new_n701), .B(new_n279), .C1(new_n221), .C2(new_n257), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n816), .B1(new_n1038), .B2(new_n1039), .C1(new_n232), .C2(new_n279), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n820), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(G107), .B2(new_n207), .C1(new_n701), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n761), .B1(new_n1042), .B2(new_n813), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1036), .B(new_n1043), .C1(new_n681), .C2(new_n1015), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n984), .A2(new_n699), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n983), .A2(new_n753), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1018), .B(new_n1044), .C1(new_n1045), .C2(new_n1046), .ZN(G393));
  NAND3_X1  g0847(.A1(new_n979), .A2(new_n981), .A3(new_n988), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n829), .B1(new_n221), .B2(new_n788), .C1(new_n839), .C2(new_n777), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n814), .B(new_n1049), .C1(G77), .C2(new_n785), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n772), .A2(new_n840), .B1(new_n781), .B2(new_n349), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n793), .A2(new_n202), .B1(new_n797), .B2(new_n259), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT109), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(KEYINPUT110), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n772), .A2(new_n1021), .B1(new_n781), .B2(new_n999), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n809), .B1(new_n778), .B2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G283), .A2(new_n997), .B1(new_n798), .B2(G294), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n285), .B(new_n807), .C1(G116), .C2(new_n785), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT110), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n768), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n813), .B1(new_n469), .B2(new_n207), .C1(new_n990), .C2(new_n242), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT108), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n761), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1066), .B(new_n1071), .C1(new_n948), .C2(new_n1015), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1048), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n986), .A2(new_n699), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n979), .A2(new_n981), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n984), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(G390));
  AOI21_X1  g0878(.A(new_n682), .B1(new_n734), .B2(new_n706), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n894), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n932), .A2(new_n925), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n924), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n751), .A2(new_n675), .A3(new_n853), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n929), .B1(new_n1084), .B2(new_n931), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n923), .B1(new_n444), .B2(new_n674), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n737), .A2(G330), .A3(new_n894), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n1085), .B2(new_n1086), .C1(new_n924), .C2(new_n1082), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n988), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n826), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n762), .B1(new_n315), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(G128), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n772), .A2(new_n1095), .B1(new_n781), .B2(new_n845), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n788), .A2(KEYINPUT53), .A3(new_n840), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT53), .B1(new_n788), .B2(new_n840), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n349), .C2(new_n843), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(G125), .C2(new_n778), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n285), .B1(new_n794), .B2(new_n202), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT115), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n793), .A2(new_n1006), .B1(new_n797), .B2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT114), .Z(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n287), .A2(new_n793), .B1(new_n781), .B2(new_n564), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n285), .B(new_n1107), .C1(G68), .C2(new_n828), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n785), .A2(G77), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n790), .A2(G87), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n797), .A2(new_n469), .B1(new_n777), .B2(new_n835), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G283), .B2(new_n831), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1094), .B1(new_n1114), .B2(new_n768), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n924), .B2(new_n765), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n853), .C1(new_n731), .C2(new_n736), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n929), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1080), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n930), .A2(new_n931), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1084), .A2(new_n931), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n928), .B1(new_n1079), .B2(new_n853), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1119), .A2(new_n1120), .B1(new_n1123), .B2(new_n1089), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n458), .A2(new_n1079), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT111), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1126), .A2(new_n915), .A3(new_n644), .A4(new_n916), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT112), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT112), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT113), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1129), .A2(new_n1131), .A3(KEYINPUT113), .A4(new_n1132), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n700), .B1(new_n1091), .B2(new_n1128), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1092), .B(new_n1116), .C1(new_n1136), .C2(new_n1139), .ZN(G378));
  NOR2_X1   g0940(.A1(new_n391), .A2(new_n672), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n405), .A2(new_n334), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n405), .B2(new_n334), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1146));
  NOR3_X1   g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n405), .A2(new_n334), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1141), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n1150), .B2(new_n1143), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n923), .A2(KEYINPUT40), .A3(new_n895), .A4(new_n894), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n906), .B1(new_n902), .B2(new_n903), .ZN(new_n1155));
  OAI211_X1 g0955(.A(G330), .B(new_n1153), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT118), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1146), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT118), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1150), .A2(new_n1143), .A3(new_n1148), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1157), .B1(new_n1156), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n908), .A2(KEYINPUT119), .A3(G330), .A4(new_n1163), .ZN(new_n1166));
  AOI221_X4 g0966(.A(new_n934), .B1(new_n1152), .B2(new_n1156), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n934), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n988), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G41), .B(new_n815), .C1(G77), .C2(new_n997), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT116), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n828), .A2(new_n314), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n795), .B2(new_n777), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n772), .A2(new_n564), .B1(new_n797), .B2(new_n264), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n469), .A2(new_n793), .B1(new_n781), .B2(new_n287), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1178), .A2(new_n1008), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1176), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT58), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n278), .B1(new_n814), .B2(new_n253), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1182), .A2(new_n1183), .B1(new_n202), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n788), .A2(new_n1103), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1186), .A2(KEYINPUT117), .B1(G150), .B2(new_n785), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(KEYINPUT117), .B2(new_n1186), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n772), .A2(new_n1189), .B1(new_n797), .B2(new_n1006), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1095), .A2(new_n781), .B1(new_n793), .B2(new_n845), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n253), .B(new_n278), .C1(new_n794), .C2(new_n349), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G124), .B2(new_n778), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT59), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1185), .B1(new_n1183), .B2(new_n1182), .C1(new_n1194), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n768), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n761), .B1(new_n202), .B2(new_n826), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n1163), .C2(new_n765), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1172), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n917), .B(new_n1126), .C1(new_n1132), .C2(new_n1124), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT57), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT57), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1205), .C1(new_n1167), .C2(new_n1171), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1204), .B1(new_n1210), .B2(new_n700), .ZN(G375));
  INV_X1    g1011(.A(new_n967), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1129), .A2(new_n1212), .A3(new_n1131), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n988), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1124), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n929), .A2(new_n764), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n762), .B1(G68), .B2(new_n1093), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G283), .A2(new_n782), .B1(new_n778), .B2(G303), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n292), .A3(new_n1005), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1033), .B(new_n1220), .C1(G97), .C2(new_n790), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n772), .A2(new_n835), .B1(new_n797), .B2(new_n287), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G116), .B2(new_n809), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT120), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT121), .Z(new_n1226));
  OAI21_X1  g1026(.A(new_n815), .B1(new_n202), .B2(new_n843), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1177), .B1(new_n1095), .B2(new_n777), .C1(new_n840), .C2(new_n797), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G159), .C2(new_n790), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n793), .A2(new_n1103), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G132), .B2(new_n831), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(new_n1006), .C2(new_n781), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1218), .B1(new_n1235), .B2(new_n768), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1216), .B1(new_n1217), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1214), .A2(new_n1237), .ZN(G381));
  OR2_X1    g1038(.A1(G375), .A2(G378), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n989), .A2(new_n1077), .A3(new_n1016), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G396), .A2(G381), .A3(G393), .A4(G384), .ZN(new_n1241));
  OR3_X1    g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(G407));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(G343), .C2(new_n1239), .ZN(G409));
  XNOR2_X1  g1043(.A(G393), .B(new_n824), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n989), .A2(new_n1016), .A3(new_n1077), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1077), .B1(new_n989), .B2(new_n1016), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(G390), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1244), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1240), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n673), .A2(G213), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n700), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1092), .A2(new_n1116), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1139), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n1135), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1254), .A2(new_n1257), .A3(new_n1203), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1127), .B1(new_n1091), .B2(new_n1128), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n934), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1169), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1260), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1203), .A2(new_n1259), .B1(new_n1212), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1172), .A2(KEYINPUT123), .A3(new_n1202), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G378), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1253), .B1(new_n1258), .B2(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1213), .B(KEYINPUT60), .Z(new_n1269));
  OAI21_X1  g1069(.A(new_n699), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1237), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G384), .B(new_n1237), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1253), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(G2897), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT62), .B1(new_n1268), .B2(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1253), .B(new_n1282), .C1(new_n1258), .C2(new_n1267), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1252), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(KEYINPUT124), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1204), .C1(new_n1210), .C2(new_n700), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1203), .A2(new_n1259), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1264), .A2(new_n1212), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1266), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1257), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1253), .A4(new_n1282), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT62), .B1(new_n1286), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1251), .B1(new_n1285), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1280), .A2(KEYINPUT126), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1278), .A2(new_n1298), .A3(new_n1279), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1268), .A2(KEYINPUT125), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1268), .A2(KEYINPUT125), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1247), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1284), .B2(KEYINPUT63), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1286), .A2(new_n1306), .A3(new_n1294), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1296), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(G378), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1275), .A2(KEYINPUT127), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1239), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1251), .A2(new_n1239), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1275), .A2(KEYINPUT127), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


