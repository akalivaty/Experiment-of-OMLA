//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  XOR2_X1   g004(.A(G127gat), .B(G134gat), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(G155gat), .B2(G162gat), .ZN(new_n210));
  AND2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n208), .A2(new_n210), .B1(KEYINPUT75), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI221_X1 g014(.A(new_n213), .B1(new_n211), .B2(KEYINPUT75), .C1(new_n208), .C2(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n207), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT4), .ZN(new_n219));
  NAND2_X1  g018(.A1(G225gat), .A2(G233gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n207), .B1(new_n222), .B2(new_n217), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n215), .A2(KEYINPUT3), .A3(new_n216), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n226));
  NAND3_X1  g025(.A1(new_n219), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n217), .A2(new_n222), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n205), .B(new_n206), .Z(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(new_n224), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n220), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT4), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n207), .A2(new_n217), .A3(KEYINPUT76), .A4(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n218), .B2(KEYINPUT4), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n215), .A2(new_n216), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n218), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n226), .B1(new_n243), .B2(new_n221), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n229), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n239), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n234), .A2(new_n236), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n225), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT78), .A3(new_n244), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n228), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G1gat), .B(G29gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT0), .ZN(new_n253));
  XNOR2_X1  g052(.A(G57gat), .B(G85gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  AOI21_X1  g054(.A(new_n203), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n251), .A2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n202), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT27), .B(G183gat), .ZN(new_n259));
  INV_X1    g058(.A(G190gat), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n259), .A2(KEYINPUT28), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G183gat), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n260), .C1(KEYINPUT68), .C2(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT26), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  OR3_X1    g080(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT25), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(KEYINPUT64), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n271), .A2(KEYINPUT25), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n297), .A3(KEYINPUT23), .ZN(new_n298));
  AND4_X1   g097(.A1(new_n288), .A2(new_n295), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n284), .B(new_n279), .C1(G183gat), .C2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n231), .B1(new_n278), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n288), .A2(new_n292), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n290), .A2(new_n289), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n305), .C1(new_n286), .C2(new_n281), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n306), .A2(KEYINPUT25), .B1(new_n300), .B2(new_n299), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n308));
  AOI21_X1  g107(.A(G190gat), .B1(new_n263), .B2(KEYINPUT68), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT28), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n276), .B(new_n275), .C1(new_n310), .C2(new_n261), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n207), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT34), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT34), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n303), .A2(new_n312), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G15gat), .B(G43gat), .Z(new_n320));
  XNOR2_X1  g119(.A(G71gat), .B(G99gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n278), .A2(new_n302), .A3(new_n231), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n207), .B1(new_n307), .B2(new_n311), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT33), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n326), .A2(KEYINPUT32), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT33), .B1(new_n313), .B2(new_n315), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n316), .B(new_n318), .C1(new_n331), .C2(new_n323), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n329), .B2(new_n332), .ZN(new_n334));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT31), .B(G50gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G22gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(new_n337), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT71), .B(G211gat), .ZN(new_n343));
  INV_X1    g142(.A(G218gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n345), .B2(KEYINPUT22), .ZN(new_n346));
  XNOR2_X1  g145(.A(G211gat), .B(G218gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(KEYINPUT72), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(KEYINPUT72), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n350), .B(new_n342), .C1(new_n345), .C2(KEYINPUT22), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n230), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n347), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n348), .B(new_n342), .C1(new_n345), .C2(KEYINPUT22), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n222), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n241), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n354), .B1(new_n359), .B2(KEYINPUT80), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n361), .A3(new_n241), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n360), .A2(new_n362), .B1(G228gat), .B2(G233gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n352), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n222), .B1(new_n365), .B2(KEYINPUT29), .ZN(new_n366));
  AOI211_X1 g165(.A(new_n364), .B(new_n354), .C1(new_n366), .C2(new_n241), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n341), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n369));
  INV_X1    g168(.A(new_n354), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n364), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n241), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n373), .A2(G228gat), .A3(G233gat), .A4(new_n370), .ZN(new_n374));
  INV_X1    g173(.A(new_n341), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n333), .A2(new_n334), .A3(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n249), .A2(KEYINPUT78), .A3(new_n244), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT78), .B1(new_n249), .B2(new_n244), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n255), .B(new_n227), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n202), .B1(new_n381), .B2(KEYINPUT79), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n227), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(new_n255), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G226gat), .ZN(new_n387));
  INV_X1    g186(.A(G233gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n307), .A2(new_n311), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n353), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n389), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n352), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n365), .B1(new_n395), .B2(new_n391), .ZN(new_n396));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT73), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(KEYINPUT30), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n396), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n400), .B(KEYINPUT74), .Z(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n402), .B1(new_n407), .B2(KEYINPUT30), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n258), .A2(new_n378), .A3(new_n386), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n381), .A2(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n385), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n413), .A2(new_n202), .B1(new_n382), .B2(new_n385), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n414), .A2(KEYINPUT83), .A3(new_n408), .A4(new_n378), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT35), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n406), .B1(new_n394), .B2(new_n396), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT30), .B1(new_n401), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(KEYINPUT30), .B2(new_n401), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n218), .A2(KEYINPUT4), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n235), .B1(new_n207), .B2(new_n217), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n232), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n221), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(KEYINPUT39), .C1(new_n221), .C2(new_n243), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT82), .A2(KEYINPUT40), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT39), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n427), .A3(new_n221), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n424), .A2(new_n255), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n220), .B1(new_n219), .B2(new_n232), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT39), .B1(new_n243), .B2(new_n221), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n255), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n257), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n377), .B1(new_n419), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n404), .A2(KEYINPUT37), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n400), .B1(new_n404), .B2(KEYINPUT37), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n406), .A2(KEYINPUT38), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n404), .B2(KEYINPUT37), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n401), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n436), .B1(new_n414), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n258), .A2(new_n386), .A3(new_n408), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n377), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n333), .A2(new_n334), .ZN(new_n448));
  NAND2_X1  g247(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OR3_X1    g252(.A1(new_n333), .A2(new_n334), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n445), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT35), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n409), .A2(new_n410), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n416), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G197gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT11), .B(G169gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  XOR2_X1   g262(.A(new_n463), .B(KEYINPUT12), .Z(new_n464));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n465), .B(KEYINPUT13), .Z(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(G1gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT16), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n471), .B2(G1gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n473), .A3(G8gat), .ZN(new_n474));
  INV_X1    g273(.A(G8gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n468), .B(new_n472), .C1(new_n469), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(G43gat), .A2(G50gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g280(.A1(G43gat), .A2(G50gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT84), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g285(.A1(G29gat), .A2(G36gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT87), .ZN(new_n488));
  AND2_X1   g287(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n489));
  NOR2_X1   g288(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n490));
  OAI22_X1  g289(.A1(new_n489), .A2(new_n490), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n492));
  INV_X1    g291(.A(G29gat), .ZN(new_n493));
  INV_X1    g292(.A(G36gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n488), .B1(new_n496), .B2(KEYINPUT86), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n486), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n484), .A2(new_n479), .A3(KEYINPUT15), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n488), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n502), .A2(new_n486), .A3(new_n496), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n478), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n506), .A2(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n507));
  INV_X1    g306(.A(new_n495), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT86), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n488), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n499), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n486), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n502), .A2(new_n486), .A3(new_n496), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(new_n477), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n466), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT89), .B(KEYINPUT17), .C1(new_n500), .C2(new_n503), .ZN(new_n518));
  OR2_X1    g317(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n519));
  NAND2_X1  g318(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n513), .A2(new_n514), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n477), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n465), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n522), .A2(new_n523), .A3(new_n505), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n517), .B1(new_n524), .B2(KEYINPUT18), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NOR4_X1   g325(.A1(new_n522), .A2(new_n505), .A3(new_n526), .A4(new_n523), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n464), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n466), .ZN(new_n529));
  INV_X1    g328(.A(new_n516), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n477), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n518), .A2(new_n521), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n478), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n465), .A3(new_n531), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n532), .B1(new_n535), .B2(new_n526), .ZN(new_n536));
  INV_X1    g335(.A(new_n464), .ZN(new_n537));
  INV_X1    g336(.A(new_n527), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n528), .A2(new_n539), .A3(KEYINPUT90), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT90), .B1(new_n528), .B2(new_n539), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n459), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(G85gat), .A3(G92gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G99gat), .B(G106gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(KEYINPUT8), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n550), .B1(new_n549), .B2(new_n554), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(new_n554), .A3(new_n550), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT95), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT96), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n549), .A2(new_n554), .ZN(new_n562));
  INV_X1    g361(.A(new_n550), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(KEYINPUT95), .A3(new_n559), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n555), .A2(new_n557), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n518), .B2(new_n521), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n570), .A2(KEYINPUT97), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n569), .A2(new_n515), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n533), .A2(KEYINPUT97), .A3(new_n561), .A4(new_n568), .ZN(new_n574));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n573), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n570), .A2(KEYINPUT97), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n577), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(KEYINPUT98), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n577), .B2(new_n580), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n594));
  INV_X1    g393(.A(G64gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(G57gat), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n596), .B(new_n598), .C1(new_n597), .C2(G64gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n602));
  NAND2_X1  g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n603), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT92), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n599), .A2(new_n604), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G57gat), .B(G64gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n603), .B(new_n601), .C1(new_n610), .C2(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n478), .B1(new_n593), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n593), .ZN(new_n614));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n613), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT93), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n617), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n565), .A2(new_n567), .B1(new_n611), .B2(new_n609), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n555), .A2(new_n556), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n627), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n634), .A2(new_n636), .A3(new_n626), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n638), .B2(new_n639), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n592), .A2(new_n625), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n544), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n414), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g454(.A(new_n475), .B1(new_n652), .B2(new_n419), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n651), .A2(new_n408), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(KEYINPUT42), .B2(new_n658), .ZN(G1325gat));
  INV_X1    g459(.A(new_n448), .ZN(new_n661));
  AOI21_X1  g460(.A(G15gat), .B1(new_n652), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n455), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT99), .Z(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n652), .B2(new_n665), .ZN(G1326gat));
  INV_X1    g465(.A(new_n377), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n459), .A2(new_n591), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n459), .A2(KEYINPUT44), .A3(new_n591), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n528), .A2(new_n539), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n648), .A2(new_n624), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n673), .A2(new_n653), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G29gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n592), .A2(new_n676), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT100), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n414), .A2(G29gat), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n459), .A2(new_n543), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT101), .ZN(G1328gat));
  NAND4_X1  g485(.A1(new_n544), .A2(new_n494), .A3(new_n419), .A4(new_n681), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(KEYINPUT102), .B2(KEYINPUT46), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n673), .A2(new_n674), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n691), .A2(new_n419), .A3(new_n677), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n494), .B2(new_n692), .ZN(G1329gat));
  NOR2_X1   g492(.A1(new_n448), .A2(G43gat), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n459), .A2(new_n543), .A3(new_n681), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT103), .Z(new_n696));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n663), .A3(new_n674), .A4(new_n677), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G43gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n698), .A3(KEYINPUT47), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1330gat));
  NAND4_X1  g502(.A1(new_n673), .A2(new_n377), .A3(new_n674), .A4(new_n677), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G50gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n667), .A2(G50gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n544), .A2(new_n681), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1331gat));
  NAND2_X1  g509(.A1(new_n528), .A2(new_n539), .ZN(new_n711));
  NOR4_X1   g510(.A1(new_n591), .A2(new_n711), .A3(new_n624), .A4(new_n648), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n459), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n414), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(new_n597), .ZN(G1332gat));
  INV_X1    g514(.A(new_n713), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n408), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT104), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n721), .B(new_n723), .ZN(G1333gat));
  NAND3_X1  g523(.A1(new_n716), .A2(G71gat), .A3(new_n663), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n713), .A2(KEYINPUT105), .A3(new_n448), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT105), .B1(new_n713), .B2(new_n448), .ZN(new_n727));
  INV_X1    g526(.A(G71gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n725), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n377), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n675), .A2(new_n624), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n647), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT107), .Z(new_n737));
  NAND2_X1  g536(.A1(new_n691), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738), .B2(new_n414), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n459), .A2(new_n591), .A3(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n459), .A2(KEYINPUT51), .A3(new_n591), .A4(new_n735), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n414), .A2(G85gat), .A3(new_n648), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT108), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n739), .B1(new_n745), .B2(new_n747), .ZN(G1336gat));
  NAND4_X1  g547(.A1(new_n673), .A2(new_n419), .A3(new_n737), .A4(new_n674), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n740), .A2(new_n752), .A3(KEYINPUT51), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n740), .B2(new_n752), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n408), .A2(G92gat), .A3(new_n648), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT52), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(new_n744), .B2(new_n755), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n750), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n750), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(G1337gat));
  OAI21_X1  g562(.A(G99gat), .B1(new_n738), .B2(new_n455), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n448), .A2(G99gat), .A3(new_n648), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n745), .B2(new_n765), .ZN(G1338gat));
  NAND4_X1  g565(.A1(new_n673), .A2(new_n377), .A3(new_n737), .A4(new_n674), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G106gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n667), .A2(G106gat), .A3(new_n648), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n753), .A2(new_n754), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n773), .A2(new_n770), .B1(G106gat), .B2(new_n767), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(new_n769), .ZN(G1339gat));
  NOR2_X1   g574(.A1(new_n649), .A2(new_n711), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n642), .B1(new_n638), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n612), .B1(new_n558), .B2(new_n560), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n612), .A2(new_n635), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT10), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n628), .B1(new_n561), .B2(new_n568), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n626), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n632), .A2(new_n637), .A3(new_n627), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n644), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n779), .A2(new_n786), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n779), .A2(new_n786), .A3(KEYINPUT55), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n525), .A2(new_n464), .A3(new_n527), .ZN(new_n795));
  INV_X1    g594(.A(new_n463), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n505), .A2(new_n516), .A3(new_n466), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n523), .B1(new_n522), .B2(new_n505), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(KEYINPUT112), .B(new_n523), .C1(new_n522), .C2(new_n505), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT113), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n463), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n539), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n591), .A2(new_n794), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n539), .A3(new_n647), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n793), .A3(new_n790), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n675), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n591), .B1(new_n811), .B2(KEYINPUT114), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n809), .C1(new_n675), .C2(new_n810), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n808), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n777), .B1(new_n815), .B2(new_n625), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n653), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n378), .A2(new_n408), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n819), .A2(G113gat), .A3(new_n675), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n816), .A2(new_n667), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n653), .A2(new_n408), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n448), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n543), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT115), .A3(G113gat), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT115), .B1(new_n824), .B2(G113gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n820), .B(new_n829), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1340gat));
  NAND2_X1  g630(.A1(new_n821), .A2(new_n823), .ZN(new_n832));
  OAI21_X1  g631(.A(G120gat), .B1(new_n832), .B2(new_n648), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n648), .A2(G120gat), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT117), .Z(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n819), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n836), .B(new_n837), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n832), .B2(new_n624), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n624), .A2(G127gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n819), .B2(new_n840), .ZN(G1342gat));
  NOR2_X1   g640(.A1(new_n592), .A2(G134gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n817), .A2(new_n818), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n832), .B2(new_n592), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n844), .A2(new_n849), .A3(new_n845), .A4(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1343gat));
  NAND2_X1  g650(.A1(new_n455), .A2(new_n377), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n419), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n817), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(G141gat), .A3(new_n542), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n663), .A2(new_n822), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n667), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n794), .B1(new_n540), .B2(new_n541), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n591), .B1(new_n860), .B2(new_n809), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n624), .B1(new_n861), .B2(new_n808), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n776), .B1(new_n862), .B2(KEYINPUT120), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT90), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n711), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n528), .A2(new_n539), .A3(KEYINPUT90), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n810), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n809), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n592), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n591), .A2(new_n794), .A3(new_n803), .A4(new_n807), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n625), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n859), .B1(new_n863), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n816), .B2(new_n377), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n856), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(new_n675), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n855), .B1(new_n877), .B2(G141gat), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n855), .A2(KEYINPUT58), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n876), .A2(new_n542), .ZN(new_n881));
  INV_X1    g680(.A(G141gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n878), .A2(new_n879), .B1(new_n880), .B2(new_n883), .ZN(G1344gat));
  OAI211_X1 g683(.A(new_n647), .B(new_n856), .C1(new_n874), .C2(new_n875), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(KEYINPUT59), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n856), .A2(new_n647), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n649), .A2(new_n543), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n377), .B1(new_n871), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n857), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n816), .A2(new_n858), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(KEYINPUT122), .B(KEYINPUT59), .C1(new_n897), .C2(new_n886), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n894), .A2(new_n857), .B1(new_n816), .B2(new_n858), .ZN(new_n900));
  OAI21_X1  g699(.A(G148gat), .B1(new_n900), .B2(new_n892), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT122), .B1(new_n901), .B2(KEYINPUT59), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n890), .B(new_n891), .C1(new_n899), .C2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n817), .A2(new_n886), .A3(new_n647), .A4(new_n853), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n876), .B2(new_n624), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n624), .A2(G155gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n854), .B2(new_n907), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n876), .B2(new_n592), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n592), .A2(G162gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n854), .B2(new_n910), .ZN(G1347gat));
  NAND2_X1  g710(.A1(new_n414), .A2(new_n419), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n448), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n821), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(G169gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(new_n542), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n816), .A2(new_n414), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n378), .A2(new_n419), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n711), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n916), .B1(new_n915), .B2(new_n921), .ZN(G1348gat));
  OAI21_X1  g721(.A(G176gat), .B1(new_n914), .B2(new_n648), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n648), .A2(G176gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n919), .B2(new_n924), .ZN(G1349gat));
  OAI21_X1  g724(.A(G183gat), .B1(new_n914), .B2(new_n624), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n917), .A2(new_n259), .A3(new_n625), .A4(new_n918), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n260), .A3(new_n591), .ZN(new_n936));
  OAI21_X1  g735(.A(G190gat), .B1(new_n914), .B2(new_n592), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n852), .A2(new_n408), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n917), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n942), .A2(G197gat), .A3(new_n675), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n895), .A2(new_n896), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n663), .A2(new_n912), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT125), .B1(new_n947), .B2(new_n542), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G197gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n947), .A2(KEYINPUT125), .A3(new_n542), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  NOR2_X1   g750(.A1(new_n648), .A2(G204gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n917), .A2(new_n941), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G204gat), .B1(new_n947), .B2(new_n648), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n625), .A3(new_n945), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n625), .A2(new_n343), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n961), .A2(new_n962), .B1(new_n942), .B2(new_n963), .ZN(G1354gat));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n344), .A3(new_n592), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n917), .A2(new_n591), .A3(new_n941), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n966), .A2(new_n344), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(G1355gat));
endmodule


