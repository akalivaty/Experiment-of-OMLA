//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n209), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n212), .B2(new_n213), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n208), .A2(new_n219), .A3(KEYINPUT87), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT87), .B1(new_n208), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT88), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(KEYINPUT88), .C1(new_n220), .C2(new_n221), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT90), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  AOI21_X1  g031(.A(G1gat), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(new_n233), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n238));
  NAND3_X1  g037(.A1(new_n224), .A2(new_n225), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n231), .B(new_n233), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n218), .B(KEYINPUT17), .C1(new_n220), .C2(new_n221), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT91), .Z(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n237), .A2(new_n242), .A3(KEYINPUT18), .A4(new_n244), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n244), .B(KEYINPUT13), .Z(new_n249));
  NOR2_X1   g048(.A1(new_n226), .A2(new_n236), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n224), .A2(new_n225), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n240), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n247), .A2(new_n259), .A3(new_n248), .A4(new_n253), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(KEYINPUT1), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(G127gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G134gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  OAI221_X1 g073(.A(new_n266), .B1(new_n267), .B2(KEYINPUT1), .C1(new_n270), .C2(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  XOR2_X1   g076(.A(G141gat), .B(G148gat), .Z(new_n278));
  INV_X1    g077(.A(G155gat), .ZN(new_n279));
  INV_X1    g078(.A(G162gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT2), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G155gat), .B(G162gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n283), .A3(new_n281), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n276), .B1(new_n277), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n286), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT79), .B1(new_n285), .B2(new_n286), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT3), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n265), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n276), .B2(new_n287), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n287), .A3(new_n293), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n276), .A2(new_n287), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n292), .B(new_n298), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n301));
  INV_X1    g100(.A(new_n276), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n289), .B2(new_n290), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n304), .B2(new_n265), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n276), .A2(new_n287), .A3(new_n293), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT4), .B1(new_n306), .B2(new_n294), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n296), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n292), .A2(new_n301), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n300), .A2(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT0), .ZN(new_n313));
  XNOR2_X1  g112(.A(G57gat), .B(G85gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  OAI21_X1  g114(.A(KEYINPUT84), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n305), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n309), .A2(new_n310), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320));
  INV_X1    g119(.A(new_n315), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n288), .A2(new_n291), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n324), .A3(new_n308), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n265), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n326), .B(KEYINPUT39), .C1(new_n265), .C2(new_n304), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT40), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT39), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n329), .A3(new_n265), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n315), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n315), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT39), .B1(new_n304), .B2(new_n265), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n265), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT40), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n323), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G169gat), .ZN(new_n338));
  INV_X1    g137(.A(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT66), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(KEYINPUT23), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n338), .A2(new_n339), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n345), .B(new_n348), .C1(new_n349), .C2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n349), .A2(KEYINPUT64), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(KEYINPUT64), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n355), .A2(new_n350), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT25), .B1(new_n343), .B2(KEYINPUT23), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n352), .A2(KEYINPUT25), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  INV_X1    g162(.A(G190gat), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n366));
  OR2_X1    g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT26), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n342), .A2(new_n368), .A3(new_n344), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n346), .B1(KEYINPUT26), .B2(new_n340), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n369), .A2(new_n370), .B1(G183gat), .B2(G190gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n361), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G197gat), .B(G204gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT73), .B(G211gat), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n381), .A2(G218gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n382), .B2(KEYINPUT22), .ZN(new_n383));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n380), .B(new_n384), .C1(new_n382), .C2(KEYINPUT22), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n378), .B(KEYINPUT76), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n379), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n386), .A2(KEYINPUT74), .A3(new_n387), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n378), .B1(new_n361), .B2(new_n373), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n389), .B1(new_n374), .B2(new_n375), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(KEYINPUT77), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n408), .B2(KEYINPUT30), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n398), .A3(KEYINPUT30), .A4(new_n402), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT85), .B1(new_n337), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n404), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n391), .A2(new_n398), .A3(new_n406), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n406), .B1(new_n391), .B2(new_n398), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n416), .A2(new_n417), .A3(new_n402), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n323), .A4(new_n336), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT3), .B1(new_n388), .B2(new_n375), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n287), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n285), .A2(new_n286), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n375), .B1(new_n427), .B2(KEYINPUT3), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n428), .A2(new_n387), .A3(new_n386), .ZN(new_n429));
  INV_X1    g228(.A(G228gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n426), .A2(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(KEYINPUT82), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n375), .C1(new_n427), .C2(KEYINPUT3), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n393), .A2(new_n433), .A3(new_n394), .A4(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n430), .A2(new_n431), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n289), .A2(new_n290), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n425), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G22gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(G22gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n432), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT31), .B(G50gat), .Z(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n444), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n443), .B1(new_n432), .B2(new_n439), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT83), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n445), .A3(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n405), .A2(KEYINPUT37), .A3(new_n407), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n403), .B1(new_n399), .B2(KEYINPUT37), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n311), .B2(new_n315), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n316), .A2(new_n462), .A3(new_n322), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n311), .A2(new_n315), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n379), .A2(new_n390), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n397), .A2(new_n396), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n466), .A2(new_n388), .B1(new_n467), .B2(new_n395), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT38), .B1(new_n468), .B2(KEYINPUT37), .ZN(new_n469));
  INV_X1    g268(.A(new_n458), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n404), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n459), .A2(new_n463), .A3(new_n465), .A4(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n414), .A2(new_n424), .A3(new_n456), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n374), .A2(new_n276), .ZN(new_n478));
  INV_X1    g277(.A(G227gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n431), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n302), .A2(new_n361), .A3(new_n373), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(KEYINPUT33), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n482), .A2(KEYINPUT32), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n481), .ZN(new_n498));
  INV_X1    g297(.A(new_n480), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n491), .B1(new_n490), .B2(new_n495), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n500), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n490), .A2(new_n495), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT34), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n505), .B2(new_n496), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n476), .B(new_n477), .C1(new_n502), .C2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n500), .B1(new_n497), .B2(new_n501), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n503), .A3(new_n496), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n474), .A4(new_n475), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n460), .B1(new_n319), .B2(new_n321), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n465), .B1(new_n512), .B2(new_n464), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n413), .A2(new_n513), .B1(new_n450), .B2(new_n454), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n473), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n413), .A2(new_n513), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n450), .A2(new_n454), .A3(new_n509), .A4(new_n508), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT35), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n422), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n463), .A2(new_n465), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n523), .B2(new_n518), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n263), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G134gat), .B(G162gat), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT101), .ZN(new_n530));
  XOR2_X1   g329(.A(G99gat), .B(G106gat), .Z(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  AND2_X1   g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n534), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT8), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n532), .B1(new_n540), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(new_n544), .B2(new_n545), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n551), .B(new_n531), .C1(new_n539), .C2(new_n538), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n550), .A2(KEYINPUT100), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT100), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n530), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT100), .ZN(new_n556));
  INV_X1    g355(.A(new_n552), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n534), .A2(new_n536), .ZN(new_n558));
  INV_X1    g357(.A(new_n537), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n531), .B1(new_n562), .B2(new_n551), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n556), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n550), .A2(KEYINPUT100), .A3(new_n552), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(KEYINPUT101), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n555), .A2(new_n241), .A3(new_n239), .A4(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n226), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n567), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n529), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT103), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(KEYINPUT103), .B(new_n529), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n570), .ZN(new_n579));
  INV_X1    g378(.A(new_n571), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n528), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n581), .A2(KEYINPUT102), .A3(new_n528), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n578), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT20), .ZN(new_n590));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  OAI221_X1 g402(.A(new_n596), .B1(new_n600), .B2(new_n601), .C1(new_n597), .C2(new_n598), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n603), .A2(KEYINPUT96), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT96), .B1(new_n603), .B2(new_n604), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n236), .B1(KEYINPUT21), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n604), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT95), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n610), .A2(new_n615), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n595), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n616), .A3(new_n594), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n431), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n569), .A2(new_n607), .A3(KEYINPUT10), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT104), .B1(new_n540), .B2(new_n549), .ZN(new_n631));
  AND4_X1   g430(.A1(new_n611), .A2(new_n631), .A3(new_n550), .A4(new_n552), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n611), .A2(new_n631), .B1(new_n550), .B2(new_n552), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n628), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n611), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n550), .A2(new_n552), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n631), .A2(new_n550), .A3(new_n611), .A4(new_n552), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n628), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT105), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n638), .A2(new_n642), .A3(new_n628), .A4(new_n639), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n626), .B1(new_n635), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT10), .B1(new_n605), .B2(new_n606), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n564), .B2(new_n565), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n638), .B2(new_n639), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n647), .A2(new_n648), .B1(new_n627), .B2(new_n431), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n649), .A2(new_n625), .A3(new_n643), .A4(new_n641), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n588), .A2(new_n622), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT106), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n588), .A2(new_n622), .A3(new_n654), .A4(new_n651), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n525), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n513), .A2(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n513), .A2(KEYINPUT107), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT109), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT108), .B(G1gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n657), .A2(new_n413), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n230), .B2(new_n665), .ZN(new_n668));
  MUX2_X1   g467(.A(new_n667), .B(new_n668), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g468(.A(new_n511), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n657), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n502), .A2(new_n506), .ZN(new_n672));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n657), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT110), .ZN(G1326gat));
  NAND3_X1  g475(.A1(new_n525), .A2(new_n455), .A3(new_n656), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n516), .A2(new_n524), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n578), .A2(new_n587), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n622), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n651), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n263), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n660), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n202), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n516), .A2(new_n524), .A3(KEYINPUT111), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n578), .A2(new_n587), .A3(KEYINPUT112), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT112), .B1(new_n578), .B2(new_n587), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n692), .A2(new_n693), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n686), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n660), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n690), .A2(new_n704), .ZN(G1328gat));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n203), .A3(new_n422), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n703), .B2(new_n413), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n210), .B1(new_n702), .B2(new_n511), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n687), .A2(new_n210), .A3(new_n672), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n516), .A2(new_n524), .A3(KEYINPUT111), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT111), .B1(new_n516), .B2(new_n524), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n715), .A3(new_n698), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n588), .B1(new_n516), .B2(new_n524), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n697), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n511), .B(new_n685), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT113), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n721), .A3(new_n511), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n720), .A2(G43gat), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n712), .A2(new_n710), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n713), .B1(new_n723), .B2(new_n724), .ZN(G1330gat));
  AOI21_X1  g524(.A(new_n211), .B1(new_n702), .B2(new_n455), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n525), .A2(new_n455), .ZN(new_n727));
  NOR4_X1   g526(.A1(new_n727), .A2(G50gat), .A3(new_n588), .A4(new_n684), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n726), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n726), .B2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1331gat));
  NAND2_X1  g532(.A1(new_n261), .A2(new_n262), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n683), .A2(new_n681), .A3(new_n734), .A4(new_n651), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n714), .A2(new_n715), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n688), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g538(.A1(new_n692), .A2(new_n693), .A3(new_n735), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT115), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n692), .A2(new_n742), .A3(new_n693), .A4(new_n735), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n422), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT49), .B(G64gat), .Z(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n692), .A2(new_n672), .A3(new_n693), .A4(new_n735), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(KEYINPUT116), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(KEYINPUT116), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n741), .A2(new_n511), .A3(new_n743), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n753), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n455), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  INV_X1    g560(.A(G85gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n622), .A2(new_n734), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n651), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n700), .B2(new_n701), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n688), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n762), .B1(new_n768), .B2(KEYINPUT117), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT117), .B2(new_n768), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n717), .B2(new_n763), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n763), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n651), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n762), .A3(new_n775), .A4(new_n688), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(G92gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n767), .B2(new_n422), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n422), .A2(new_n778), .A3(new_n775), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n772), .B2(new_n773), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n779), .A2(KEYINPUT52), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1337gat));
  INV_X1    g583(.A(G99gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n774), .A2(new_n785), .A3(new_n672), .A4(new_n775), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n767), .A2(new_n511), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n785), .ZN(G1338gat));
  NOR3_X1   g587(.A1(new_n456), .A2(G106gat), .A3(new_n651), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n456), .B(new_n766), .C1(new_n700), .C2(new_n701), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT119), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n455), .B(new_n765), .C1(new_n716), .C2(new_n718), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n790), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n797), .A2(new_n800), .A3(new_n790), .A4(new_n791), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n795), .A2(new_n799), .A3(new_n801), .ZN(G1339gat));
  NOR2_X1   g601(.A1(new_n652), .A2(new_n734), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n625), .B1(new_n635), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n629), .A2(new_n634), .A3(new_n628), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n649), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT55), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n650), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n250), .A2(new_n252), .A3(new_n249), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n244), .B1(new_n237), .B2(new_n242), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n258), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n262), .A2(new_n815), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n812), .A2(new_n263), .B1(new_n651), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n694), .B2(new_n695), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n681), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n578), .A2(new_n587), .A3(KEYINPUT112), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n812), .A2(new_n816), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n803), .B1(new_n824), .B2(new_n683), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n518), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n660), .A2(new_n422), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n263), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT120), .B(G113gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n829), .B(new_n830), .ZN(G1340gat));
  NOR2_X1   g630(.A1(new_n828), .A2(new_n651), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g632(.A1(new_n828), .A2(new_n683), .ZN(new_n834));
  NOR2_X1   g633(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(G1342gat));
  NAND3_X1  g635(.A1(new_n826), .A2(new_n681), .A3(new_n827), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(G134gat), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT56), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(G134gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1343gat));
  OR3_X1    g640(.A1(new_n825), .A2(KEYINPUT122), .A3(new_n660), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT122), .B1(new_n825), .B2(new_n660), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n670), .A2(new_n455), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n422), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n263), .A2(G141gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n670), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n825), .B2(new_n456), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n455), .A2(KEYINPUT57), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n817), .A2(new_n588), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n622), .B1(new_n823), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n803), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n849), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n734), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n847), .A2(new_n848), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  XOR2_X1   g658(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n860));
  XNOR2_X1  g659(.A(new_n859), .B(new_n860), .ZN(G1344gat));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  INV_X1    g662(.A(new_n849), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n811), .A2(new_n650), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT55), .B1(new_n805), .B2(new_n807), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n262), .A3(new_n815), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n854), .B1(new_n588), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n683), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n653), .A2(new_n263), .A3(new_n655), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n455), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n825), .A2(new_n852), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n775), .B(new_n864), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n863), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n651), .B(new_n849), .C1(new_n851), .C2(new_n856), .ZN(new_n878));
  INV_X1    g677(.A(G148gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT59), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n694), .A2(new_n868), .A3(new_n695), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n816), .A2(new_n651), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n867), .B2(new_n734), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n820), .B2(new_n821), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n683), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n803), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n455), .ZN(new_n890));
  INV_X1    g689(.A(new_n856), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n775), .B(new_n864), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(KEYINPUT124), .A3(new_n880), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n876), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n846), .A2(G148gat), .A3(new_n651), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n862), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n875), .A2(G148gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT59), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n877), .B(new_n881), .C1(new_n857), .C2(new_n775), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT124), .B1(new_n892), .B2(new_n880), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n895), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(KEYINPUT125), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n896), .A2(new_n903), .ZN(G1345gat));
  NAND3_X1  g703(.A1(new_n847), .A2(new_n279), .A3(new_n622), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n857), .A2(new_n622), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n279), .B2(new_n906), .ZN(G1346gat));
  NAND3_X1  g706(.A1(new_n847), .A2(new_n280), .A3(new_n681), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n857), .A2(new_n696), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n280), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n688), .A2(new_n413), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n826), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n263), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(new_n338), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n651), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(new_n339), .ZN(G1349gat));
  INV_X1    g715(.A(new_n912), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n622), .ZN(new_n918));
  INV_X1    g717(.A(G183gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n363), .B2(new_n918), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n912), .B2(new_n588), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT61), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n364), .A3(new_n696), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1351gat));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n670), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n872), .A2(new_n455), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n850), .ZN(new_n931));
  INV_X1    g730(.A(new_n874), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n928), .B1(new_n934), .B2(new_n263), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(KEYINPUT126), .A3(new_n734), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(G197gat), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n844), .A2(new_n688), .A3(new_n413), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n889), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n263), .A2(G197gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  OR3_X1    g740(.A1(new_n939), .A2(G204gat), .A3(new_n651), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  OAI21_X1  g742(.A(G204gat), .B1(new_n934), .B2(new_n651), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1353gat));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n932), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  INV_X1    g747(.A(new_n929), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n622), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n933), .B2(new_n622), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n622), .A3(new_n949), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n950), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OR3_X1    g756(.A1(new_n939), .A2(new_n381), .A3(new_n683), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n934), .B2(new_n588), .ZN(new_n960));
  INV_X1    g759(.A(G218gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n696), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n939), .B2(new_n962), .ZN(G1355gat));
endmodule


