

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780;

  XNOR2_X1 U371 ( .A(n550), .B(KEYINPUT39), .ZN(n552) );
  NAND2_X4 U372 ( .A1(n645), .A2(G953), .ZN(n667) );
  XNOR2_X2 U373 ( .A(n663), .B(n664), .ZN(n665) );
  XNOR2_X2 U374 ( .A(n373), .B(n641), .ZN(n643) );
  XNOR2_X2 U375 ( .A(n656), .B(n655), .ZN(n657) );
  AND2_X2 U376 ( .A1(n591), .A2(n410), .ZN(n363) );
  NAND2_X1 U377 ( .A1(n418), .A2(n421), .ZN(n417) );
  XNOR2_X1 U378 ( .A(n627), .B(n626), .ZN(n421) );
  AND2_X2 U379 ( .A1(n368), .A2(n545), .ZN(n549) );
  XOR2_X2 U380 ( .A(KEYINPUT80), .B(n588), .Z(n589) );
  XNOR2_X2 U381 ( .A(n516), .B(n770), .ZN(n651) );
  XNOR2_X2 U382 ( .A(n615), .B(KEYINPUT1), .ZN(n413) );
  OR2_X2 U383 ( .A1(n675), .A2(G902), .ZN(n543) );
  NOR2_X1 U384 ( .A1(n727), .A2(n575), .ZN(n613) );
  NOR2_X1 U385 ( .A1(n593), .A2(n733), .ZN(n597) );
  INV_X1 U386 ( .A(G953), .ZN(n773) );
  XNOR2_X1 U387 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n348) );
  AND2_X1 U388 ( .A1(n351), .A2(n378), .ZN(n349) );
  AND2_X1 U389 ( .A1(n364), .A2(n592), .ZN(n350) );
  AND2_X2 U390 ( .A1(n389), .A2(n680), .ZN(n388) );
  NAND2_X2 U391 ( .A1(n419), .A2(n417), .ZN(n416) );
  XNOR2_X2 U392 ( .A(n617), .B(KEYINPUT110), .ZN(n690) );
  NOR2_X2 U393 ( .A1(n748), .A2(G953), .ZN(n749) );
  XNOR2_X2 U394 ( .A(n622), .B(KEYINPUT41), .ZN(n722) );
  AND2_X2 U395 ( .A1(n712), .A2(n370), .ZN(n622) );
  NAND2_X2 U396 ( .A1(n405), .A2(n404), .ZN(n607) );
  XNOR2_X2 U397 ( .A(n570), .B(n367), .ZN(n582) );
  AND2_X1 U398 ( .A1(n621), .A2(n360), .ZN(n628) );
  INV_X1 U399 ( .A(n609), .ZN(n351) );
  INV_X1 U400 ( .A(n724), .ZN(n596) );
  NAND2_X1 U401 ( .A1(n727), .A2(n726), .ZN(n723) );
  NAND2_X1 U402 ( .A1(n362), .A2(n352), .ZN(n415) );
  XNOR2_X1 U403 ( .A(n597), .B(n359), .ZN(n372) );
  NOR2_X1 U404 ( .A1(n593), .A2(n599), .ZN(n600) );
  NAND2_X1 U405 ( .A1(n351), .A2(n382), .ZN(n429) );
  NOR2_X1 U406 ( .A1(n722), .A2(n690), .ZN(n624) );
  INV_X1 U407 ( .A(KEYINPUT22), .ZN(n367) );
  INV_X1 U408 ( .A(KEYINPUT47), .ZN(n361) );
  INV_X1 U409 ( .A(n628), .ZN(n362) );
  AND2_X1 U410 ( .A1(n628), .A2(n629), .ZN(n418) );
  NOR2_X1 U411 ( .A1(n601), .A2(n716), .ZN(n603) );
  NOR2_X1 U412 ( .A1(n631), .A2(n630), .ZN(n632) );
  AND2_X1 U413 ( .A1(n427), .A2(n428), .ZN(n621) );
  AND2_X1 U414 ( .A1(n392), .A2(n548), .ZN(n630) );
  NOR2_X1 U415 ( .A1(n372), .A2(n600), .ZN(n601) );
  AND2_X1 U416 ( .A1(n429), .A2(n424), .ZN(n427) );
  AND2_X1 U417 ( .A1(n399), .A2(n400), .ZN(n394) );
  XNOR2_X1 U418 ( .A(n620), .B(n361), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n624), .B(n623), .ZN(n406) );
  NAND2_X1 U420 ( .A1(n549), .A2(n712), .ZN(n550) );
  NAND2_X1 U421 ( .A1(n712), .A2(n404), .ZN(n371) );
  AND2_X1 U422 ( .A1(n724), .A2(n571), .ZN(n572) );
  XNOR2_X1 U423 ( .A(n369), .B(n348), .ZN(n368) );
  AND2_X1 U424 ( .A1(n544), .A2(n615), .ZN(n545) );
  NAND2_X1 U425 ( .A1(n730), .A2(n404), .ZN(n369) );
  BUF_X1 U426 ( .A(n730), .Z(n396) );
  XNOR2_X1 U427 ( .A(n492), .B(n481), .ZN(n758) );
  XNOR2_X1 U428 ( .A(n353), .B(n480), .ZN(n492) );
  XNOR2_X1 U429 ( .A(n354), .B(KEYINPUT3), .ZN(n353) );
  INV_X1 U430 ( .A(n629), .ZN(n352) );
  XNOR2_X1 U431 ( .A(G134), .B(G131), .ZN(n768) );
  XNOR2_X1 U432 ( .A(G140), .B(G131), .ZN(n446) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n454) );
  XNOR2_X1 U434 ( .A(G110), .B(G107), .ZN(n479) );
  INV_X1 U435 ( .A(KEYINPUT31), .ZN(n359) );
  NAND2_X1 U436 ( .A1(n582), .A2(n383), .ZN(n358) );
  XNOR2_X2 U437 ( .A(G113), .B(KEYINPUT93), .ZN(n354) );
  XNOR2_X1 U438 ( .A(n540), .B(n355), .ZN(n662) );
  XNOR2_X1 U439 ( .A(n758), .B(n356), .ZN(n355) );
  XNOR2_X1 U440 ( .A(n357), .B(n379), .ZN(n356) );
  XNOR2_X1 U441 ( .A(n483), .B(n484), .ZN(n357) );
  XNOR2_X2 U442 ( .A(n493), .B(n445), .ZN(n540) );
  XNOR2_X2 U443 ( .A(n765), .B(n478), .ZN(n493) );
  XNOR2_X2 U444 ( .A(n477), .B(KEYINPUT4), .ZN(n765) );
  XNOR2_X2 U445 ( .A(n358), .B(KEYINPUT32), .ZN(n410) );
  NAND2_X1 U446 ( .A1(n625), .A2(n406), .ZN(n627) );
  XNOR2_X2 U447 ( .A(n555), .B(n554), .ZN(n625) );
  NOR2_X1 U448 ( .A1(n690), .A2(n716), .ZN(n619) );
  NAND2_X1 U449 ( .A1(n388), .A2(n390), .ZN(n387) );
  NAND2_X1 U450 ( .A1(n350), .A2(n363), .ZN(n391) );
  AND2_X2 U451 ( .A1(n364), .A2(n591), .ZN(n411) );
  XNOR2_X1 U452 ( .A(n364), .B(G122), .ZN(G24) );
  XNOR2_X2 U453 ( .A(n402), .B(n590), .ZN(n364) );
  XNOR2_X2 U454 ( .A(n365), .B(n385), .ZN(n742) );
  NAND2_X1 U455 ( .A1(n366), .A2(n413), .ZN(n365) );
  AND2_X2 U456 ( .A1(n586), .A2(n585), .ZN(n366) );
  XNOR2_X2 U457 ( .A(n574), .B(n573), .ZN(n586) );
  XNOR2_X2 U458 ( .A(n543), .B(n542), .ZN(n615) );
  NAND2_X1 U459 ( .A1(n582), .A2(n572), .ZN(n591) );
  XNOR2_X1 U460 ( .A(n410), .B(G119), .ZN(G21) );
  NOR2_X1 U461 ( .A1(n714), .A2(n556), .ZN(n370) );
  NOR2_X1 U462 ( .A1(n716), .A2(n371), .ZN(n717) );
  BUF_X1 U463 ( .A(n642), .Z(n373) );
  XNOR2_X2 U464 ( .A(n637), .B(KEYINPUT75), .ZN(n710) );
  NAND2_X1 U465 ( .A1(n618), .A2(n563), .ZN(n374) );
  NAND2_X1 U466 ( .A1(n618), .A2(n563), .ZN(n564) );
  XNOR2_X1 U467 ( .A(n374), .B(KEYINPUT0), .ZN(n375) );
  BUF_X1 U468 ( .A(n586), .Z(n376) );
  INV_X1 U469 ( .A(n377), .ZN(n593) );
  XNOR2_X1 U470 ( .A(n374), .B(n433), .ZN(n377) );
  XNOR2_X1 U471 ( .A(n564), .B(n433), .ZN(n569) );
  XNOR2_X2 U472 ( .A(n607), .B(n558), .ZN(n618) );
  XNOR2_X1 U473 ( .A(G119), .B(G116), .ZN(n480) );
  INV_X1 U474 ( .A(KEYINPUT66), .ZN(n441) );
  AND2_X1 U475 ( .A1(n633), .A2(KEYINPUT66), .ZN(n443) );
  NAND2_X1 U476 ( .A1(n634), .A2(n439), .ZN(n438) );
  NAND2_X1 U477 ( .A1(KEYINPUT2), .A2(n441), .ZN(n439) );
  INV_X1 U478 ( .A(n416), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n576) );
  XNOR2_X1 U480 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U481 ( .A(G128), .B(G119), .ZN(n509) );
  INV_X1 U482 ( .A(KEYINPUT65), .ZN(n639) );
  XOR2_X1 U483 ( .A(G122), .B(G104), .Z(n447) );
  XNOR2_X1 U484 ( .A(G125), .B(G146), .ZN(n486) );
  XOR2_X1 U485 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n484) );
  NAND2_X1 U486 ( .A1(n586), .A2(n613), .ZN(n423) );
  INV_X1 U487 ( .A(KEYINPUT106), .ZN(n422) );
  INV_X1 U488 ( .A(G128), .ZN(n468) );
  XOR2_X1 U489 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n452) );
  XNOR2_X1 U490 ( .A(KEYINPUT16), .B(G122), .ZN(n481) );
  XNOR2_X1 U491 ( .A(G116), .B(G134), .ZN(n462) );
  XOR2_X1 U492 ( .A(G107), .B(G122), .Z(n463) );
  NAND2_X1 U493 ( .A1(n634), .A2(n441), .ZN(n435) );
  AND2_X1 U494 ( .A1(n442), .A2(n437), .ZN(n436) );
  NAND2_X1 U495 ( .A1(n440), .A2(n438), .ZN(n437) );
  NAND2_X1 U496 ( .A1(n518), .A2(n441), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n635), .B(KEYINPUT85), .ZN(n636) );
  NAND2_X1 U498 ( .A1(n408), .A2(n407), .ZN(n635) );
  XNOR2_X1 U499 ( .A(n511), .B(n510), .ZN(n514) );
  NOR2_X1 U500 ( .A1(n608), .A2(n611), .ZN(n430) );
  NAND2_X1 U501 ( .A1(n351), .A2(n431), .ZN(n426) );
  NAND2_X1 U502 ( .A1(n431), .A2(n432), .ZN(n425) );
  INV_X1 U503 ( .A(KEYINPUT28), .ZN(n395) );
  NAND2_X1 U504 ( .A1(n605), .A2(n727), .ZN(n680) );
  XNOR2_X1 U505 ( .A(n578), .B(n577), .ZN(n609) );
  INV_X1 U506 ( .A(n413), .ZN(n724) );
  INV_X1 U507 ( .A(n556), .ZN(n404) );
  NOR2_X1 U508 ( .A1(n596), .A2(n556), .ZN(n378) );
  XOR2_X1 U509 ( .A(n486), .B(n485), .Z(n379) );
  AND2_X1 U510 ( .A1(n568), .A2(n726), .ZN(n380) );
  AND2_X1 U511 ( .A1(n582), .A2(n581), .ZN(n381) );
  AND2_X1 U512 ( .A1(n430), .A2(n596), .ZN(n382) );
  NOR2_X1 U513 ( .A1(n584), .A2(n376), .ZN(n383) );
  AND2_X1 U514 ( .A1(n596), .A2(n425), .ZN(n384) );
  XNOR2_X1 U515 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n385) );
  XOR2_X1 U516 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n386) );
  INV_X1 U517 ( .A(n518), .ZN(n634) );
  XNOR2_X2 U518 ( .A(n387), .B(KEYINPUT45), .ZN(n701) );
  NAND2_X1 U519 ( .A1(n409), .A2(n412), .ZN(n389) );
  AND2_X2 U520 ( .A1(n391), .A2(n606), .ZN(n390) );
  OR2_X1 U521 ( .A1(n444), .A2(n435), .ZN(n434) );
  NOR2_X1 U522 ( .A1(n414), .A2(n633), .ZN(n407) );
  NAND2_X1 U523 ( .A1(n420), .A2(n352), .ZN(n419) );
  NAND2_X1 U524 ( .A1(n552), .A2(n694), .ZN(n555) );
  BUF_X1 U525 ( .A(n742), .Z(n393) );
  INV_X1 U526 ( .A(n592), .ZN(n412) );
  XNOR2_X1 U527 ( .A(n614), .B(n395), .ZN(n616) );
  NOR2_X2 U528 ( .A1(n416), .A2(n414), .ZN(n772) );
  XNOR2_X1 U529 ( .A(n349), .B(n386), .ZN(n392) );
  NAND2_X1 U530 ( .A1(n426), .A2(n384), .ZN(n428) );
  NAND2_X1 U531 ( .A1(n394), .A2(n397), .ZN(n403) );
  NAND2_X1 U532 ( .A1(n632), .A2(n415), .ZN(n414) );
  NAND2_X1 U533 ( .A1(n398), .A2(n377), .ZN(n397) );
  NOR2_X1 U534 ( .A1(n742), .A2(n401), .ZN(n398) );
  NAND2_X1 U535 ( .A1(n742), .A2(n401), .ZN(n399) );
  NAND2_X1 U536 ( .A1(n375), .A2(n401), .ZN(n400) );
  INV_X1 U537 ( .A(KEYINPUT34), .ZN(n401) );
  NAND2_X1 U538 ( .A1(n403), .A2(n589), .ZN(n402) );
  INV_X1 U539 ( .A(n557), .ZN(n405) );
  XNOR2_X1 U540 ( .A(n491), .B(n490), .ZN(n557) );
  XNOR2_X1 U541 ( .A(n406), .B(G137), .ZN(G39) );
  NAND2_X1 U542 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U543 ( .A(n421), .ZN(n420) );
  XNOR2_X1 U544 ( .A(n502), .B(n501), .ZN(n642) );
  XNOR2_X2 U545 ( .A(n503), .B(G472), .ZN(n574) );
  INV_X1 U546 ( .A(n612), .ZN(n424) );
  NAND2_X1 U547 ( .A1(n428), .A2(n429), .ZN(n698) );
  NAND2_X1 U548 ( .A1(n608), .A2(n611), .ZN(n431) );
  INV_X1 U549 ( .A(n611), .ZN(n432) );
  INV_X1 U550 ( .A(KEYINPUT0), .ZN(n433) );
  NAND2_X1 U551 ( .A1(n701), .A2(n772), .ZN(n444) );
  NAND2_X1 U552 ( .A1(n444), .A2(n443), .ZN(n442) );
  NAND2_X1 U553 ( .A1(n436), .A2(n434), .ZN(n638) );
  NOR2_X1 U554 ( .A1(n662), .A2(n634), .ZN(n491) );
  XOR2_X1 U555 ( .A(n756), .B(KEYINPUT70), .Z(n445) );
  INV_X1 U556 ( .A(KEYINPUT46), .ZN(n626) );
  INV_X1 U557 ( .A(G110), .ZN(n508) );
  INV_X1 U558 ( .A(KEYINPUT107), .ZN(n577) );
  INV_X1 U559 ( .A(n376), .ZN(n581) );
  XNOR2_X1 U560 ( .A(n493), .B(n494), .ZN(n502) );
  BUF_X1 U561 ( .A(n618), .Z(n692) );
  XNOR2_X1 U562 ( .A(n486), .B(KEYINPUT10), .ZN(n515) );
  XNOR2_X1 U563 ( .A(n447), .B(n446), .ZN(n449) );
  NOR2_X1 U564 ( .A1(G953), .A2(G237), .ZN(n496) );
  NAND2_X1 U565 ( .A1(G214), .A2(n496), .ZN(n448) );
  XNOR2_X1 U566 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U567 ( .A(n515), .B(n450), .Z(n457) );
  XNOR2_X1 U568 ( .A(KEYINPUT101), .B(KEYINPUT12), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U570 ( .A(n453), .B(KEYINPUT102), .Z(n455) );
  XNOR2_X1 U571 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n457), .B(n456), .ZN(n656) );
  NOR2_X1 U573 ( .A1(G902), .A2(n656), .ZN(n459) );
  XNOR2_X1 U574 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n458) );
  XNOR2_X1 U575 ( .A(n459), .B(n458), .ZN(n461) );
  INV_X1 U576 ( .A(G475), .ZN(n460) );
  XNOR2_X1 U577 ( .A(n461), .B(n460), .ZN(n567) );
  INV_X1 U578 ( .A(n567), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n463), .B(n462), .ZN(n467) );
  XOR2_X1 U580 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n465) );
  XNOR2_X1 U581 ( .A(KEYINPUT9), .B(KEYINPUT105), .ZN(n464) );
  XNOR2_X1 U582 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U583 ( .A(n467), .B(n466), .Z(n473) );
  XNOR2_X2 U584 ( .A(G143), .B(KEYINPUT64), .ZN(n469) );
  XNOR2_X2 U585 ( .A(n469), .B(n468), .ZN(n477) );
  NAND2_X1 U586 ( .A1(G234), .A2(n773), .ZN(n470) );
  XOR2_X1 U587 ( .A(KEYINPUT8), .B(n470), .Z(n512) );
  NAND2_X1 U588 ( .A1(G217), .A2(n512), .ZN(n471) );
  XNOR2_X1 U589 ( .A(n477), .B(n471), .ZN(n472) );
  XNOR2_X1 U590 ( .A(n473), .B(n472), .ZN(n649) );
  INV_X1 U591 ( .A(G902), .ZN(n517) );
  NAND2_X1 U592 ( .A1(n649), .A2(n517), .ZN(n475) );
  INV_X1 U593 ( .A(G478), .ZN(n474) );
  XNOR2_X1 U594 ( .A(n475), .B(n474), .ZN(n565) );
  NOR2_X1 U595 ( .A1(n476), .A2(n565), .ZN(n587) );
  XNOR2_X1 U596 ( .A(KEYINPUT67), .B(G101), .ZN(n478) );
  XNOR2_X1 U597 ( .A(n479), .B(G104), .ZN(n756) );
  NAND2_X1 U598 ( .A1(G224), .A2(n773), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n482), .B(KEYINPUT78), .ZN(n483) );
  XNOR2_X1 U600 ( .A(KEYINPUT90), .B(KEYINPUT94), .ZN(n485) );
  XNOR2_X1 U601 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n487) );
  XNOR2_X1 U602 ( .A(n487), .B(G902), .ZN(n518) );
  NOR2_X1 U603 ( .A1(G902), .A2(G237), .ZN(n488) );
  XNOR2_X1 U604 ( .A(n488), .B(KEYINPUT72), .ZN(n504) );
  INV_X1 U605 ( .A(G210), .ZN(n489) );
  NOR2_X1 U606 ( .A1(n504), .A2(n489), .ZN(n490) );
  BUF_X1 U607 ( .A(n557), .Z(n548) );
  INV_X1 U608 ( .A(n548), .ZN(n579) );
  NAND2_X1 U609 ( .A1(n587), .A2(n579), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n492), .B(G137), .ZN(n494) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(KEYINPUT99), .ZN(n495) );
  XNOR2_X1 U612 ( .A(n768), .B(G146), .ZN(n538) );
  XNOR2_X1 U613 ( .A(n495), .B(n538), .ZN(n500) );
  XOR2_X1 U614 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n498) );
  NAND2_X1 U615 ( .A1(G210), .A2(n496), .ZN(n497) );
  XNOR2_X1 U616 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U617 ( .A(n500), .B(n499), .Z(n501) );
  NAND2_X1 U618 ( .A1(n642), .A2(n517), .ZN(n503) );
  BUF_X2 U619 ( .A(n574), .Z(n730) );
  INV_X1 U620 ( .A(n504), .ZN(n505) );
  AND2_X1 U621 ( .A1(n505), .A2(G214), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT97), .B(KEYINPUT23), .Z(n507) );
  XNOR2_X1 U623 ( .A(KEYINPUT77), .B(KEYINPUT24), .ZN(n506) );
  XNOR2_X1 U624 ( .A(n507), .B(n506), .ZN(n511) );
  NAND2_X1 U625 ( .A1(n512), .A2(G221), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n514), .B(n513), .ZN(n516) );
  INV_X1 U627 ( .A(G140), .ZN(n580) );
  XNOR2_X1 U628 ( .A(n580), .B(G137), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n515), .B(n534), .ZN(n770) );
  NAND2_X1 U630 ( .A1(n651), .A2(n517), .ZN(n523) );
  NAND2_X1 U631 ( .A1(G234), .A2(n518), .ZN(n519) );
  XNOR2_X1 U632 ( .A(KEYINPUT20), .B(n519), .ZN(n524) );
  NAND2_X1 U633 ( .A1(G217), .A2(n524), .ZN(n521) );
  INV_X1 U634 ( .A(KEYINPUT25), .ZN(n520) );
  XNOR2_X1 U635 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X2 U636 ( .A(n523), .B(n522), .ZN(n727) );
  INV_X1 U637 ( .A(n727), .ZN(n583) );
  NAND2_X1 U638 ( .A1(n524), .A2(G221), .ZN(n527) );
  INV_X1 U639 ( .A(KEYINPUT98), .ZN(n525) );
  XNOR2_X1 U640 ( .A(n525), .B(KEYINPUT21), .ZN(n526) );
  XNOR2_X1 U641 ( .A(n527), .B(n526), .ZN(n726) );
  NAND2_X1 U642 ( .A1(G237), .A2(G234), .ZN(n528) );
  XNOR2_X1 U643 ( .A(n528), .B(KEYINPUT14), .ZN(n529) );
  NAND2_X1 U644 ( .A1(G952), .A2(n529), .ZN(n741) );
  NOR2_X1 U645 ( .A1(G953), .A2(n741), .ZN(n561) );
  AND2_X1 U646 ( .A1(G953), .A2(n529), .ZN(n530) );
  NAND2_X1 U647 ( .A1(G902), .A2(n530), .ZN(n559) );
  NOR2_X1 U648 ( .A1(G900), .A2(n559), .ZN(n531) );
  NOR2_X1 U649 ( .A1(n561), .A2(n531), .ZN(n532) );
  XNOR2_X1 U650 ( .A(n532), .B(KEYINPUT81), .ZN(n533) );
  NAND2_X1 U651 ( .A1(n726), .A2(n533), .ZN(n575) );
  NOR2_X1 U652 ( .A1(n583), .A2(n575), .ZN(n544) );
  INV_X1 U653 ( .A(n534), .ZN(n536) );
  NAND2_X1 U654 ( .A1(n773), .A2(G227), .ZN(n535) );
  XNOR2_X1 U655 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U656 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U657 ( .A(n540), .B(n539), .ZN(n675) );
  INV_X1 U658 ( .A(KEYINPUT69), .ZN(n541) );
  XNOR2_X1 U659 ( .A(n541), .B(G469), .ZN(n542) );
  INV_X1 U660 ( .A(n549), .ZN(n546) );
  NOR2_X1 U661 ( .A1(n547), .A2(n546), .ZN(n612) );
  XOR2_X1 U662 ( .A(G143), .B(n612), .Z(G45) );
  XNOR2_X2 U663 ( .A(n548), .B(KEYINPUT38), .ZN(n712) );
  INV_X1 U664 ( .A(n552), .ZN(n551) );
  OR2_X1 U665 ( .A1(n567), .A2(n565), .ZN(n685) );
  NOR2_X1 U666 ( .A1(n551), .A2(n685), .ZN(n631) );
  XOR2_X1 U667 ( .A(G134), .B(n631), .Z(G36) );
  AND2_X1 U668 ( .A1(n567), .A2(n565), .ZN(n694) );
  XOR2_X1 U669 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n553) );
  XNOR2_X1 U670 ( .A(n553), .B(KEYINPUT111), .ZN(n554) );
  XNOR2_X1 U671 ( .A(n625), .B(G131), .ZN(G33) );
  XNOR2_X1 U672 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n558) );
  XOR2_X1 U673 ( .A(G898), .B(KEYINPUT95), .Z(n759) );
  NOR2_X1 U674 ( .A1(n559), .A2(n759), .ZN(n560) );
  OR2_X1 U675 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U676 ( .A(n562), .B(KEYINPUT96), .ZN(n563) );
  INV_X1 U677 ( .A(n565), .ZN(n566) );
  OR2_X1 U678 ( .A1(n567), .A2(n566), .ZN(n714) );
  INV_X1 U679 ( .A(n714), .ZN(n568) );
  NAND2_X1 U680 ( .A1(n569), .A2(n380), .ZN(n570) );
  NOR2_X1 U681 ( .A1(n396), .A2(n727), .ZN(n571) );
  XNOR2_X1 U682 ( .A(n591), .B(G110), .ZN(G12) );
  INV_X1 U683 ( .A(KEYINPUT6), .ZN(n573) );
  NAND2_X1 U684 ( .A1(n576), .A2(n694), .ZN(n578) );
  XNOR2_X1 U685 ( .A(n630), .B(n580), .ZN(G42) );
  NAND2_X1 U686 ( .A1(n596), .A2(n583), .ZN(n584) );
  INV_X1 U687 ( .A(n723), .ZN(n585) );
  INV_X1 U688 ( .A(n587), .ZN(n588) );
  XNOR2_X1 U689 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n590) );
  NOR2_X1 U690 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n592) );
  INV_X1 U691 ( .A(n396), .ZN(n594) );
  NOR2_X1 U692 ( .A1(n594), .A2(n723), .ZN(n595) );
  NAND2_X1 U693 ( .A1(n596), .A2(n595), .ZN(n733) );
  NOR2_X1 U694 ( .A1(n396), .A2(n723), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n598), .A2(n615), .ZN(n599) );
  INV_X1 U696 ( .A(n694), .ZN(n689) );
  AND2_X1 U697 ( .A1(n689), .A2(n685), .ZN(n716) );
  AND2_X1 U698 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n602) );
  NOR2_X1 U699 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U700 ( .A1(n381), .A2(n724), .ZN(n604) );
  XNOR2_X1 U701 ( .A(n604), .B(KEYINPUT87), .ZN(n605) );
  BUF_X1 U702 ( .A(n607), .Z(n608) );
  XNOR2_X1 U703 ( .A(KEYINPUT88), .B(KEYINPUT114), .ZN(n610) );
  XOR2_X1 U704 ( .A(n610), .B(KEYINPUT36), .Z(n611) );
  NAND2_X1 U705 ( .A1(n730), .A2(n613), .ZN(n614) );
  NAND2_X1 U706 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U707 ( .A1(n619), .A2(n692), .ZN(n620) );
  XNOR2_X1 U708 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n623) );
  XOR2_X1 U709 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n629) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n636), .A2(n701), .ZN(n637) );
  NOR2_X2 U712 ( .A1(n638), .A2(n710), .ZN(n640) );
  XNOR2_X2 U713 ( .A(n640), .B(n639), .ZN(n672) );
  NAND2_X1 U714 ( .A1(n672), .A2(G472), .ZN(n644) );
  XOR2_X1 U715 ( .A(KEYINPUT91), .B(KEYINPUT62), .Z(n641) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n646) );
  INV_X1 U717 ( .A(G952), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n646), .A2(n667), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U720 ( .A1(n672), .A2(G478), .ZN(n648) );
  XOR2_X1 U721 ( .A(n649), .B(n648), .Z(n650) );
  INV_X1 U722 ( .A(n667), .ZN(n678) );
  NOR2_X1 U723 ( .A1(n650), .A2(n678), .ZN(G63) );
  NAND2_X1 U724 ( .A1(n672), .A2(G217), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n653), .A2(n667), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n654), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U728 ( .A1(n672), .A2(G475), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n655) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n659), .A2(n667), .ZN(n661) );
  XOR2_X1 U732 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(G60) );
  NAND2_X1 U734 ( .A1(n672), .A2(G210), .ZN(n666) );
  BUF_X1 U735 ( .A(n662), .Z(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n671) );
  XNOR2_X1 U739 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n669) );
  XOR2_X1 U740 ( .A(n669), .B(KEYINPUT86), .Z(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G51) );
  BUF_X1 U742 ( .A(n672), .Z(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(G469), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(G54) );
  XNOR2_X1 U748 ( .A(G101), .B(n680), .ZN(G3) );
  NAND2_X1 U749 ( .A1(n600), .A2(n694), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(G104), .ZN(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n683) );
  INV_X1 U752 ( .A(n685), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n600), .A2(n696), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(G107), .B(n684), .ZN(G9) );
  NOR2_X1 U756 ( .A1(n690), .A2(n685), .ZN(n686) );
  AND2_X1 U757 ( .A1(n686), .A2(n692), .ZN(n687) );
  XNOR2_X1 U758 ( .A(G128), .B(n687), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT29), .ZN(G30) );
  NOR2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  AND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U762 ( .A(G146), .B(n693), .Z(G48) );
  NAND2_X1 U763 ( .A1(n372), .A2(n694), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(G113), .ZN(G15) );
  NAND2_X1 U765 ( .A1(n372), .A2(n696), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(G116), .ZN(G18) );
  XOR2_X1 U767 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n700) );
  XNOR2_X1 U768 ( .A(n698), .B(G125), .ZN(n699) );
  XNOR2_X1 U769 ( .A(n700), .B(n699), .ZN(G27) );
  INV_X1 U770 ( .A(n772), .ZN(n703) );
  BUF_X2 U771 ( .A(n701), .Z(n750) );
  NOR2_X1 U772 ( .A1(n750), .A2(KEYINPUT83), .ZN(n702) );
  NOR2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U774 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n705) );
  OR2_X1 U775 ( .A1(n704), .A2(n705), .ZN(n708) );
  OR2_X1 U776 ( .A1(n750), .A2(n705), .ZN(n706) );
  NAND2_X1 U777 ( .A1(n706), .A2(KEYINPUT83), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U780 ( .A(KEYINPUT84), .B(n711), .Z(n747) );
  NOR2_X1 U781 ( .A1(n712), .A2(n404), .ZN(n713) );
  NOR2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U783 ( .A(n715), .B(KEYINPUT116), .ZN(n718) );
  NOR2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U785 ( .A(KEYINPUT117), .B(n719), .Z(n720) );
  NOR2_X1 U786 ( .A1(n720), .A2(n393), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n721), .B(KEYINPUT118), .ZN(n738) );
  NAND2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U789 ( .A(n725), .B(KEYINPUT50), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U791 ( .A(KEYINPUT49), .B(n728), .Z(n729) );
  NOR2_X1 U792 ( .A1(n396), .A2(n729), .ZN(n731) );
  NAND2_X1 U793 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U794 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U795 ( .A(KEYINPUT51), .B(n735), .ZN(n736) );
  NOR2_X1 U796 ( .A1(n722), .A2(n736), .ZN(n737) );
  NOR2_X1 U797 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U798 ( .A(n739), .B(KEYINPUT52), .ZN(n740) );
  NOR2_X1 U799 ( .A1(n741), .A2(n740), .ZN(n745) );
  NOR2_X1 U800 ( .A1(n722), .A2(n393), .ZN(n743) );
  XOR2_X1 U801 ( .A(KEYINPUT119), .B(n743), .Z(n744) );
  NOR2_X1 U802 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U803 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n749), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U805 ( .A1(n750), .A2(n773), .ZN(n754) );
  NAND2_X1 U806 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U807 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U808 ( .A1(n752), .A2(n759), .ZN(n753) );
  NAND2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U810 ( .A(n755), .B(KEYINPUT125), .ZN(n764) );
  XOR2_X1 U811 ( .A(G101), .B(n756), .Z(n757) );
  XNOR2_X1 U812 ( .A(n758), .B(n757), .ZN(n761) );
  NOR2_X1 U813 ( .A1(n759), .A2(n773), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U815 ( .A(n762), .B(KEYINPUT124), .Z(n763) );
  XNOR2_X1 U816 ( .A(n764), .B(n763), .ZN(G69) );
  BUF_X1 U817 ( .A(n765), .Z(n766) );
  INV_X1 U818 ( .A(KEYINPUT126), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U820 ( .A(n766), .B(n769), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n775) );
  XOR2_X1 U822 ( .A(n775), .B(n772), .Z(n774) );
  NAND2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n780) );
  XNOR2_X1 U824 ( .A(G227), .B(n775), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(G953), .ZN(n778) );
  XOR2_X1 U827 ( .A(KEYINPUT127), .B(n778), .Z(n779) );
  NAND2_X1 U828 ( .A1(n780), .A2(n779), .ZN(G72) );
endmodule

