

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U554 ( .A1(n718), .A2(n717), .ZN(n762) );
  OR2_X1 U555 ( .A1(n730), .A2(n729), .ZN(n739) );
  XNOR2_X1 U556 ( .A(n719), .B(KEYINPUT96), .ZN(n720) );
  INV_X2 U557 ( .A(n762), .ZN(n747) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n539), .ZN(n868) );
  NOR2_X2 U559 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  INV_X1 U560 ( .A(KEYINPUT99), .ZN(n740) );
  NOR2_X1 U561 ( .A1(n619), .A2(n524), .ZN(n640) );
  XNOR2_X1 U562 ( .A(n741), .B(n740), .ZN(n745) );
  XNOR2_X1 U563 ( .A(KEYINPUT72), .B(KEYINPUT13), .ZN(n559) );
  NOR2_X1 U564 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U565 ( .A(n560), .B(n559), .ZN(n564) );
  NOR2_X1 U566 ( .A1(G651), .A2(n619), .ZN(n637) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n644) );
  AND2_X1 U568 ( .A1(n538), .A2(n537), .ZN(n684) );
  NOR2_X2 U569 ( .A1(n566), .A2(n565), .ZN(n927) );
  NAND2_X1 U570 ( .A1(n644), .A2(G89), .ZN(n520) );
  XNOR2_X1 U571 ( .A(n520), .B(KEYINPUT4), .ZN(n522) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n619) );
  INV_X1 U573 ( .A(G651), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G76), .A2(n640), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U576 ( .A(n523), .B(KEYINPUT5), .ZN(n530) );
  NOR2_X1 U577 ( .A1(G543), .A2(n524), .ZN(n525) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n525), .Z(n636) );
  NAND2_X1 U579 ( .A1(G63), .A2(n636), .ZN(n527) );
  NAND2_X1 U580 ( .A1(G51), .A2(n637), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U582 ( .A(KEYINPUT6), .B(n528), .Z(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U584 ( .A(n531), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U585 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X2 U586 ( .A(KEYINPUT17), .B(n532), .Z(n869) );
  NAND2_X1 U587 ( .A1(G137), .A2(n869), .ZN(n534) );
  INV_X1 U588 ( .A(G2104), .ZN(n539) );
  INV_X1 U589 ( .A(G2105), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n539), .A2(n536), .ZN(n864) );
  NAND2_X1 U591 ( .A1(G113), .A2(n864), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U593 ( .A(n535), .B(KEYINPUT65), .ZN(n538) );
  NOR2_X1 U594 ( .A1(G2104), .A2(n536), .ZN(n865) );
  NAND2_X1 U595 ( .A1(G125), .A2(n865), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G101), .A2(n868), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n540), .B(KEYINPUT64), .ZN(n541) );
  XOR2_X1 U598 ( .A(n541), .B(KEYINPUT23), .Z(n683) );
  AND2_X1 U599 ( .A1(n684), .A2(n683), .ZN(G160) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U601 ( .A1(G123), .A2(n865), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n542), .B(KEYINPUT18), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G111), .A2(n864), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n543), .B(KEYINPUT78), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n868), .A2(G99), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G135), .A2(n869), .ZN(n546) );
  XNOR2_X1 U608 ( .A(KEYINPUT77), .B(n546), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n999) );
  XNOR2_X1 U611 ( .A(G2096), .B(n999), .ZN(n551) );
  OR2_X1 U612 ( .A1(G2100), .A2(n551), .ZN(G156) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U618 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n554) );
  INV_X1 U619 ( .A(G223), .ZN(n821) );
  NAND2_X1 U620 ( .A1(G567), .A2(n821), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G234) );
  NAND2_X1 U622 ( .A1(n637), .A2(G43), .ZN(n555) );
  XNOR2_X1 U623 ( .A(KEYINPUT73), .B(n555), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n644), .A2(G81), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n556), .B(KEYINPUT12), .ZN(n558) );
  NAND2_X1 U626 ( .A1(G68), .A2(n640), .ZN(n557) );
  NAND2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(KEYINPUT71), .Z(n562) );
  NAND2_X1 U629 ( .A1(G56), .A2(n636), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n927), .A2(G860), .ZN(G153) );
  NAND2_X1 U633 ( .A1(G64), .A2(n636), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G52), .A2(n637), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G77), .A2(n640), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G90), .A2(n644), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT67), .B(n574), .ZN(G301) );
  NAND2_X1 U642 ( .A1(G301), .A2(G868), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT74), .ZN(n585) );
  INV_X1 U644 ( .A(G868), .ZN(n655) );
  NAND2_X1 U645 ( .A1(n637), .A2(G54), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G79), .A2(n640), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G92), .A2(n644), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G66), .A2(n636), .ZN(n578) );
  XNOR2_X1 U650 ( .A(KEYINPUT75), .B(n578), .ZN(n579) );
  NOR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT15), .B(n583), .Z(n914) );
  NAND2_X1 U654 ( .A1(n655), .A2(n914), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U656 ( .A(KEYINPUT76), .B(n586), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G65), .A2(n636), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT68), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G78), .A2(n640), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G91), .A2(n644), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G53), .A2(n637), .ZN(n590) );
  XNOR2_X1 U663 ( .A(KEYINPUT69), .B(n590), .ZN(n591) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(G299) );
  NOR2_X1 U666 ( .A1(G286), .A2(n655), .ZN(n596) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(G297) );
  INV_X1 U669 ( .A(G860), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n597), .A2(G559), .ZN(n598) );
  INV_X1 U671 ( .A(n914), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n598), .A2(n603), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U674 ( .A1(n603), .A2(G868), .ZN(n600) );
  NOR2_X1 U675 ( .A1(G559), .A2(n600), .ZN(n602) );
  AND2_X1 U676 ( .A1(n655), .A2(n927), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G282) );
  XOR2_X1 U678 ( .A(n927), .B(KEYINPUT79), .Z(n605) );
  NAND2_X1 U679 ( .A1(G559), .A2(n603), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n605), .B(n604), .ZN(n653) );
  XOR2_X1 U681 ( .A(n653), .B(KEYINPUT80), .Z(n606) );
  NOR2_X1 U682 ( .A1(G860), .A2(n606), .ZN(n614) );
  NAND2_X1 U683 ( .A1(G67), .A2(n636), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G55), .A2(n637), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G93), .A2(n644), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT81), .B(n609), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n640), .A2(G80), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n656) );
  XOR2_X1 U691 ( .A(n614), .B(n656), .Z(G145) );
  NAND2_X1 U692 ( .A1(G49), .A2(n637), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U695 ( .A(KEYINPUT82), .B(n617), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n636), .A2(n618), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n619), .A2(G87), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(G288) );
  NAND2_X1 U699 ( .A1(G73), .A2(n640), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT2), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G61), .A2(n636), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G86), .A2(n644), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G48), .A2(n637), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT83), .B(n625), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G75), .A2(n640), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G88), .A2(n644), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G62), .A2(n636), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G50), .A2(n637), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G60), .A2(n636), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G47), .A2(n637), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G72), .A2(n640), .ZN(n641) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(n641), .Z(n642) );
  NOR2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n644), .A2(G85), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(G290) );
  XOR2_X1 U723 ( .A(G299), .B(G305), .Z(n647) );
  XNOR2_X1 U724 ( .A(G288), .B(n647), .ZN(n648) );
  XOR2_X1 U725 ( .A(n648), .B(KEYINPUT19), .Z(n650) );
  XNOR2_X1 U726 ( .A(G166), .B(KEYINPUT84), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(G290), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n652), .B(n656), .ZN(n889) );
  XOR2_X1 U730 ( .A(n889), .B(n653), .Z(n654) );
  NOR2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n658) );
  NOR2_X1 U732 ( .A1(G868), .A2(n656), .ZN(n657) );
  NOR2_X1 U733 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2084), .A2(G2078), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n660), .ZN(n662) );
  XOR2_X1 U737 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U739 ( .A1(G2072), .A2(n663), .ZN(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U741 ( .A1(G220), .A2(G219), .ZN(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT22), .B(n664), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n665), .A2(G96), .ZN(n666) );
  NOR2_X1 U744 ( .A1(G218), .A2(n666), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT86), .B(n667), .Z(n827) );
  NAND2_X1 U746 ( .A1(n827), .A2(G2106), .ZN(n671) );
  NAND2_X1 U747 ( .A1(G120), .A2(G108), .ZN(n668) );
  NOR2_X1 U748 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(G69), .A2(n669), .ZN(n826) );
  NAND2_X1 U750 ( .A1(G567), .A2(n826), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT87), .B(n672), .ZN(G319) );
  INV_X1 U753 ( .A(G319), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n673) );
  XNOR2_X1 U755 ( .A(KEYINPUT88), .B(n673), .ZN(n674) );
  NOR2_X1 U756 ( .A1(n675), .A2(n674), .ZN(n825) );
  NAND2_X1 U757 ( .A1(n825), .A2(G36), .ZN(n676) );
  XOR2_X1 U758 ( .A(KEYINPUT89), .B(n676), .Z(G176) );
  NAND2_X1 U759 ( .A1(G102), .A2(n868), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G138), .A2(n869), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G114), .A2(n864), .ZN(n680) );
  NAND2_X1 U763 ( .A1(G126), .A2(n865), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U765 ( .A1(n682), .A2(n681), .ZN(G164) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  INV_X1 U767 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U768 ( .A(G1986), .B(G290), .ZN(n926) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n718) );
  AND2_X1 U770 ( .A1(G40), .A2(n683), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n716) );
  NOR2_X1 U772 ( .A1(n718), .A2(n716), .ZN(n816) );
  NAND2_X1 U773 ( .A1(n926), .A2(n816), .ZN(n805) );
  NAND2_X1 U774 ( .A1(G104), .A2(n868), .ZN(n687) );
  NAND2_X1 U775 ( .A1(G140), .A2(n869), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U777 ( .A(KEYINPUT34), .B(n688), .ZN(n694) );
  NAND2_X1 U778 ( .A1(G116), .A2(n864), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G128), .A2(n865), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U781 ( .A(KEYINPUT90), .B(n691), .Z(n692) );
  XNOR2_X1 U782 ( .A(KEYINPUT35), .B(n692), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U784 ( .A(n695), .B(KEYINPUT36), .Z(n696) );
  XNOR2_X1 U785 ( .A(KEYINPUT91), .B(n696), .ZN(n877) );
  XNOR2_X1 U786 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  NOR2_X1 U787 ( .A1(n877), .A2(n814), .ZN(n1008) );
  NAND2_X1 U788 ( .A1(n816), .A2(n1008), .ZN(n697) );
  XNOR2_X1 U789 ( .A(KEYINPUT92), .B(n697), .ZN(n812) );
  NAND2_X1 U790 ( .A1(G95), .A2(n868), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G131), .A2(n869), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U793 ( .A(KEYINPUT93), .B(n700), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G107), .A2(n864), .ZN(n702) );
  NAND2_X1 U795 ( .A1(G119), .A2(n865), .ZN(n701) );
  AND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n878) );
  AND2_X1 U798 ( .A1(n878), .A2(G1991), .ZN(n713) );
  NAND2_X1 U799 ( .A1(G117), .A2(n864), .ZN(n706) );
  NAND2_X1 U800 ( .A1(G129), .A2(n865), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n868), .A2(G105), .ZN(n707) );
  XOR2_X1 U803 ( .A(KEYINPUT38), .B(n707), .Z(n708) );
  NOR2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n869), .A2(G141), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n882) );
  AND2_X1 U807 ( .A1(n882), .A2(G1996), .ZN(n712) );
  NOR2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n990) );
  INV_X1 U809 ( .A(n816), .ZN(n714) );
  NOR2_X1 U810 ( .A1(n990), .A2(n714), .ZN(n808) );
  INV_X1 U811 ( .A(n808), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n812), .A2(n715), .ZN(n803) );
  INV_X1 U813 ( .A(n716), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n747), .A2(G1996), .ZN(n719) );
  XNOR2_X1 U815 ( .A(n720), .B(KEYINPUT26), .ZN(n725) );
  NAND2_X1 U816 ( .A1(G2067), .A2(n747), .ZN(n721) );
  XNOR2_X1 U817 ( .A(n721), .B(KEYINPUT98), .ZN(n723) );
  NAND2_X1 U818 ( .A1(G1348), .A2(n762), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n735), .A2(n914), .ZN(n724) );
  NAND2_X1 U821 ( .A1(n725), .A2(n724), .ZN(n730) );
  INV_X1 U822 ( .A(n927), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n762), .A2(G1341), .ZN(n726) );
  XNOR2_X1 U824 ( .A(n726), .B(KEYINPUT97), .ZN(n727) );
  OR2_X1 U825 ( .A1(n728), .A2(n727), .ZN(n729) );
  INV_X1 U826 ( .A(G2072), .ZN(n967) );
  NOR2_X1 U827 ( .A1(n762), .A2(n967), .ZN(n732) );
  XOR2_X1 U828 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n731) );
  XNOR2_X1 U829 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U830 ( .A1(n762), .A2(G1956), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G299), .A2(n742), .ZN(n737) );
  NOR2_X1 U833 ( .A1(n735), .A2(n914), .ZN(n736) );
  NOR2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U836 ( .A1(G299), .A2(n742), .ZN(n743) );
  XNOR2_X1 U837 ( .A(KEYINPUT28), .B(n743), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U839 ( .A(n746), .B(KEYINPUT29), .ZN(n751) );
  OR2_X1 U840 ( .A1(n747), .A2(G1961), .ZN(n749) );
  XNOR2_X1 U841 ( .A(KEYINPUT25), .B(G2078), .ZN(n973) );
  NAND2_X1 U842 ( .A1(n747), .A2(n973), .ZN(n748) );
  NAND2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n753) );
  AND2_X1 U844 ( .A1(G171), .A2(n753), .ZN(n750) );
  NOR2_X1 U845 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U846 ( .A(n752), .B(KEYINPUT100), .ZN(n761) );
  NOR2_X1 U847 ( .A1(G171), .A2(n753), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G8), .A2(n762), .ZN(n799) );
  NOR2_X1 U849 ( .A1(G1966), .A2(n799), .ZN(n772) );
  NOR2_X1 U850 ( .A1(G2084), .A2(n762), .ZN(n770) );
  NOR2_X1 U851 ( .A1(n772), .A2(n770), .ZN(n754) );
  NAND2_X1 U852 ( .A1(G8), .A2(n754), .ZN(n755) );
  XNOR2_X1 U853 ( .A(KEYINPUT30), .B(n755), .ZN(n756) );
  NOR2_X1 U854 ( .A1(G168), .A2(n756), .ZN(n757) );
  NOR2_X1 U855 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U856 ( .A(KEYINPUT31), .B(n759), .ZN(n760) );
  OR2_X2 U857 ( .A1(n761), .A2(n760), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n774), .A2(G286), .ZN(n767) );
  NOR2_X1 U859 ( .A1(G1971), .A2(n799), .ZN(n764) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U861 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U862 ( .A1(n765), .A2(G303), .ZN(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n768), .A2(G8), .ZN(n769) );
  XNOR2_X1 U865 ( .A(n769), .B(KEYINPUT32), .ZN(n777) );
  AND2_X1 U866 ( .A1(G8), .A2(n770), .ZN(n771) );
  NOR2_X1 U867 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U868 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U869 ( .A(KEYINPUT101), .B(n775), .Z(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n792) );
  NOR2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n924) );
  NOR2_X1 U872 ( .A1(G1971), .A2(G303), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n924), .A2(n778), .ZN(n780) );
  INV_X1 U874 ( .A(KEYINPUT33), .ZN(n779) );
  AND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n792), .A2(n781), .ZN(n785) );
  INV_X1 U877 ( .A(n799), .ZN(n782) );
  NAND2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n917) );
  AND2_X1 U879 ( .A1(n782), .A2(n917), .ZN(n783) );
  OR2_X1 U880 ( .A1(KEYINPUT33), .A2(n783), .ZN(n784) );
  NAND2_X1 U881 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n924), .A2(KEYINPUT33), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n786), .A2(n799), .ZN(n787) );
  NOR2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U885 ( .A(G1981), .B(G305), .Z(n911) );
  NAND2_X1 U886 ( .A1(n789), .A2(n911), .ZN(n795) );
  NOR2_X1 U887 ( .A1(G2090), .A2(G303), .ZN(n790) );
  NAND2_X1 U888 ( .A1(G8), .A2(n790), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n793), .A2(n799), .ZN(n794) );
  NAND2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n801) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U893 ( .A(n796), .B(KEYINPUT94), .Z(n797) );
  XNOR2_X1 U894 ( .A(KEYINPUT24), .B(n797), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n819) );
  XNOR2_X1 U898 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n811) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n882), .ZN(n1004) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n878), .ZN(n998) );
  NOR2_X1 U902 ( .A1(n806), .A2(n998), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n1004), .A2(n809), .ZN(n810) );
  XNOR2_X1 U905 ( .A(n811), .B(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n877), .A2(n814), .ZN(n1006) );
  NAND2_X1 U908 ( .A1(n815), .A2(n1006), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U911 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n823) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(n823), .Z(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U918 ( .A(G108), .B(KEYINPUT111), .ZN(G238) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(G2678), .Z(n829) );
  XNOR2_X1 U925 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT42), .B(G2090), .Z(n831) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U930 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2096), .B(G2100), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U933 ( .A(G2084), .B(G2078), .Z(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1956), .B(G1961), .Z(n839) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n849) );
  XOR2_X1 U938 ( .A(KEYINPUT108), .B(KEYINPUT110), .Z(n841) );
  XNOR2_X1 U939 ( .A(G1991), .B(KEYINPUT41), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U941 ( .A(G1976), .B(G1981), .Z(n843) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1971), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U944 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT109), .B(G2474), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U948 ( .A1(G124), .A2(n865), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U950 ( .A1(n864), .A2(G112), .ZN(n851) );
  NAND2_X1 U951 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U952 ( .A1(G100), .A2(n868), .ZN(n854) );
  NAND2_X1 U953 ( .A1(G136), .A2(n869), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U955 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U956 ( .A1(G103), .A2(n868), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G139), .A2(n869), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G115), .A2(n864), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G127), .A2(n865), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n992) );
  NAND2_X1 U964 ( .A1(G118), .A2(n864), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G130), .A2(n865), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G106), .A2(n868), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G142), .A2(n869), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n875), .B(n999), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n992), .B(n876), .ZN(n881) );
  XNOR2_X1 U974 ( .A(G160), .B(n877), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U976 ( .A(n881), .B(n880), .ZN(n887) );
  XOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  XOR2_X1 U978 ( .A(n882), .B(G162), .Z(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U980 ( .A(G164), .B(n885), .Z(n886) );
  XNOR2_X1 U981 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U982 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U983 ( .A(n914), .B(n889), .ZN(n891) );
  XNOR2_X1 U984 ( .A(G171), .B(n927), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U986 ( .A(G286), .B(n892), .Z(n893) );
  NOR2_X1 U987 ( .A1(G37), .A2(n893), .ZN(G397) );
  XNOR2_X1 U988 ( .A(G2451), .B(G2427), .ZN(n903) );
  XOR2_X1 U989 ( .A(KEYINPUT103), .B(G2443), .Z(n895) );
  XNOR2_X1 U990 ( .A(G2435), .B(G2438), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U992 ( .A(G2454), .B(G2430), .Z(n897) );
  XNOR2_X1 U993 ( .A(G1341), .B(G1348), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U996 ( .A(G2446), .B(KEYINPUT104), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  NAND2_X1 U999 ( .A1(n904), .A2(G14), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n910), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  INV_X1 U1008 ( .A(n910), .ZN(G401) );
  XOR2_X1 U1009 ( .A(KEYINPUT56), .B(G16), .Z(n935) );
  XNOR2_X1 U1010 ( .A(G1966), .B(G168), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n913), .B(KEYINPUT57), .ZN(n923) );
  XNOR2_X1 U1013 ( .A(n914), .B(G1348), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(G299), .B(G1956), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1017 ( .A(G1961), .B(G171), .Z(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT116), .B(n919), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n933) );
  XOR2_X1 U1021 ( .A(n924), .B(KEYINPUT117), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n931) );
  XOR2_X1 U1023 ( .A(n927), .B(G1341), .Z(n929) );
  XNOR2_X1 U1024 ( .A(G303), .B(G1971), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n1020) );
  XNOR2_X1 U1029 ( .A(G1986), .B(KEYINPUT124), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(n936), .B(G24), .ZN(n942) );
  XNOR2_X1 U1031 ( .A(G1976), .B(KEYINPUT122), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(G23), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G22), .B(G1971), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(KEYINPUT123), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(KEYINPUT58), .B(n943), .ZN(n961) );
  XNOR2_X1 U1038 ( .A(KEYINPUT119), .B(G1981), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n944), .B(G6), .ZN(n949) );
  XOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .Z(n945) );
  XNOR2_X1 U1041 ( .A(G4), .B(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(G19), .B(G1341), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G20), .B(G1956), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(KEYINPUT118), .B(n950), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(n953), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(KEYINPUT60), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G5), .B(G1961), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT121), .B(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n962), .B(KEYINPUT125), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n963) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n965), .ZN(n989) );
  XOR2_X1 U1060 ( .A(G2067), .B(G26), .Z(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(G28), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT114), .B(n967), .Z(n968) );
  XNOR2_X1 U1063 ( .A(G33), .B(n968), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G1991), .B(G25), .Z(n972) );
  XOR2_X1 U1066 ( .A(G1996), .B(G32), .Z(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G27), .B(n973), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(KEYINPUT53), .ZN(n981) );
  XOR2_X1 U1072 ( .A(G2084), .B(G34), .Z(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT54), .B(n979), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G35), .B(G2090), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT55), .B(n984), .Z(n985) );
  NOR2_X1 U1078 ( .A1(G29), .A2(n985), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT115), .B(n986), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(G11), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n1018) );
  XNOR2_X1 U1082 ( .A(G160), .B(G2084), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n1002) );
  XNOR2_X1 U1084 ( .A(G164), .B(G2078), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G2072), .B(n992), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT112), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT50), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1011) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n1005), .Z(n1007) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT113), .B(n1013), .ZN(n1015) );
  INV_X1 U1100 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1021), .Z(n1022) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

