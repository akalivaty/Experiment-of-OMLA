

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G2105), .A2(n527), .ZN(n528) );
  BUF_X1 U556 ( .A(n1007), .Z(n521) );
  XNOR2_X1 U557 ( .A(n528), .B(KEYINPUT66), .ZN(n1007) );
  NOR2_X1 U558 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U559 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X2 U560 ( .A1(n582), .A2(n581), .ZN(G164) );
  NOR2_X2 U561 ( .A1(n532), .A2(n531), .ZN(n1003) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n747) );
  XNOR2_X1 U563 ( .A(n748), .B(n747), .ZN(n753) );
  NAND2_X1 U564 ( .A1(n716), .A2(n715), .ZN(n754) );
  BUF_X1 U565 ( .A(n754), .Z(n766) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  NOR2_X1 U567 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U568 ( .A1(G651), .A2(n626), .ZN(n651) );
  NOR2_X1 U569 ( .A1(n536), .A2(n535), .ZN(G160) );
  XNOR2_X1 U570 ( .A(n522), .B(KEYINPUT67), .ZN(n523) );
  XNOR2_X2 U571 ( .A(n523), .B(KEYINPUT17), .ZN(n1006) );
  NAND2_X1 U572 ( .A1(G137), .A2(n1006), .ZN(n525) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n1002) );
  NAND2_X1 U574 ( .A1(G113), .A2(n1002), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U576 ( .A(n526), .B(KEYINPUT68), .ZN(n536) );
  INV_X1 U577 ( .A(KEYINPUT23), .ZN(n530) );
  XNOR2_X1 U578 ( .A(KEYINPUT65), .B(G2104), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n1007), .A2(G101), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n530), .B(n529), .ZN(n534) );
  INV_X1 U581 ( .A(G2105), .ZN(n532) );
  XOR2_X1 U582 ( .A(G2104), .B(KEYINPUT65), .Z(n531) );
  NAND2_X1 U583 ( .A1(G125), .A2(n1003), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X1 U585 ( .A(G651), .ZN(n546) );
  NOR2_X1 U586 ( .A1(G543), .A2(n546), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n537), .Z(n650) );
  NAND2_X1 U588 ( .A1(n650), .A2(G63), .ZN(n538) );
  XNOR2_X1 U589 ( .A(KEYINPUT77), .B(n538), .ZN(n541) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NAND2_X1 U591 ( .A1(n651), .A2(G51), .ZN(n539) );
  XOR2_X1 U592 ( .A(n539), .B(KEYINPUT78), .Z(n540) );
  NOR2_X1 U593 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U594 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  XNOR2_X1 U595 ( .A(n543), .B(KEYINPUT79), .ZN(n551) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U597 ( .A1(G89), .A2(n646), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n544), .B(KEYINPUT76), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT4), .ZN(n548) );
  NOR2_X1 U600 ( .A1(n626), .A2(n546), .ZN(n647) );
  NAND2_X1 U601 ( .A1(G76), .A2(n647), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U603 ( .A(KEYINPUT5), .B(n549), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U605 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G64), .A2(n650), .ZN(n554) );
  NAND2_X1 U608 ( .A1(G52), .A2(n651), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G90), .A2(n646), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G77), .A2(n647), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U614 ( .A1(n559), .A2(n558), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n1003), .A2(G123), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n560), .B(KEYINPUT18), .ZN(n567) );
  NAND2_X1 U617 ( .A1(G135), .A2(n1006), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G99), .A2(n521), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G111), .A2(n1002), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT81), .B(n563), .ZN(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n1013) );
  XNOR2_X1 U624 ( .A(G2096), .B(n1013), .ZN(n568) );
  OR2_X1 U625 ( .A1(G2100), .A2(n568), .ZN(G156) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(G65), .A2(n650), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G53), .A2(n651), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G91), .A2(n646), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G78), .A2(n647), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n743) );
  INV_X1 U636 ( .A(n743), .ZN(G299) );
  NAND2_X1 U637 ( .A1(G138), .A2(n1006), .ZN(n575) );
  XNOR2_X1 U638 ( .A(n575), .B(KEYINPUT90), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n1003), .A2(G126), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT89), .B(n576), .Z(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n1002), .A2(G114), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n521), .A2(G102), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G94), .A2(G452), .ZN(n583) );
  XOR2_X1 U646 ( .A(KEYINPUT70), .B(n583), .Z(G173) );
  XOR2_X1 U647 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n585) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G223) );
  INV_X1 U650 ( .A(G223), .ZN(n827) );
  NAND2_X1 U651 ( .A1(n827), .A2(G567), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  NAND2_X1 U653 ( .A1(n650), .A2(G56), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n587), .Z(n593) );
  NAND2_X1 U655 ( .A1(n646), .A2(G81), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G68), .A2(n647), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n591), .Z(n592) );
  NOR2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n594), .B(KEYINPUT72), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G43), .A2(n651), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n1023) );
  INV_X1 U664 ( .A(G860), .ZN(n611) );
  OR2_X1 U665 ( .A1(n1023), .A2(n611), .ZN(G153) );
  NAND2_X1 U666 ( .A1(G92), .A2(n646), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G79), .A2(n647), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G66), .A2(n650), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G54), .A2(n651), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n604) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(KEYINPUT15), .B(n605), .ZN(n841) );
  NOR2_X1 U676 ( .A1(G868), .A2(n841), .ZN(n607) );
  INV_X1 U677 ( .A(G868), .ZN(n657) );
  NOR2_X1 U678 ( .A1(G171), .A2(n657), .ZN(n606) );
  NOR2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT75), .B(n608), .ZN(G284) );
  NOR2_X1 U681 ( .A1(G286), .A2(n657), .ZN(n610) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n612), .A2(n841), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT80), .ZN(n614) );
  XNOR2_X1 U687 ( .A(KEYINPUT16), .B(n614), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n1023), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n841), .A2(G868), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G559), .A2(n615), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G61), .A2(n650), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G86), .A2(n646), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n647), .A2(G73), .ZN(n620) );
  XOR2_X1 U696 ( .A(KEYINPUT2), .B(n620), .Z(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U698 ( .A(KEYINPUT83), .B(n623), .Z(n625) );
  NAND2_X1 U699 ( .A1(n651), .A2(G48), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(G305) );
  NAND2_X1 U701 ( .A1(G49), .A2(n651), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G87), .A2(n626), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n650), .A2(n629), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G651), .A2(G74), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G62), .A2(n650), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G88), .A2(n646), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n647), .A2(G75), .ZN(n634) );
  XOR2_X1 U711 ( .A(KEYINPUT84), .B(n634), .Z(n635) );
  NOR2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n651), .A2(G50), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(G303) );
  INV_X1 U715 ( .A(G303), .ZN(G166) );
  NAND2_X1 U716 ( .A1(G60), .A2(n650), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G47), .A2(n651), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U719 ( .A(KEYINPUT69), .B(n641), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G85), .A2(n646), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G72), .A2(n647), .ZN(n642) );
  AND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U724 ( .A1(G93), .A2(n646), .ZN(n649) );
  NAND2_X1 U725 ( .A1(G80), .A2(n647), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n649), .A2(n648), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G67), .A2(n650), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G55), .A2(n651), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U731 ( .A(KEYINPUT82), .B(n656), .Z(n960) );
  NAND2_X1 U732 ( .A1(n657), .A2(n960), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(KEYINPUT86), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n660) );
  XNOR2_X1 U735 ( .A(G288), .B(n960), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U737 ( .A(G305), .B(n661), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n743), .B(G166), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(G290), .ZN(n1019) );
  NAND2_X1 U741 ( .A1(n841), .A2(G559), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(n1023), .ZN(n958) );
  XNOR2_X1 U743 ( .A(n1019), .B(n958), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT87), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(KEYINPUT20), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U756 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(G96), .A2(n676), .ZN(n961) );
  NAND2_X1 U758 ( .A1(n961), .A2(G2106), .ZN(n680) );
  NAND2_X1 U759 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U760 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G108), .A2(n678), .ZN(n962) );
  NAND2_X1 U762 ( .A1(n962), .A2(G567), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n680), .A2(n679), .ZN(n1032) );
  NOR2_X1 U764 ( .A1(n681), .A2(n1032), .ZN(n682) );
  XNOR2_X1 U765 ( .A(n682), .B(KEYINPUT88), .ZN(n830) );
  NAND2_X1 U766 ( .A1(G36), .A2(n830), .ZN(G176) );
  XNOR2_X1 U767 ( .A(G1986), .B(G290), .ZN(n858) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n822) );
  NAND2_X1 U771 ( .A1(n858), .A2(n822), .ZN(n810) );
  NAND2_X1 U772 ( .A1(G131), .A2(n1006), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G95), .A2(n521), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n1002), .A2(G107), .ZN(n687) );
  NAND2_X1 U776 ( .A1(G119), .A2(n1003), .ZN(n686) );
  NAND2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n998) );
  INV_X1 U779 ( .A(G1991), .ZN(n866) );
  NOR2_X1 U780 ( .A1(n998), .A2(n866), .ZN(n701) );
  NAND2_X1 U781 ( .A1(n521), .A2(G105), .ZN(n692) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(KEYINPUT93), .Z(n690) );
  XNOR2_X1 U783 ( .A(KEYINPUT92), .B(n690), .ZN(n691) );
  XNOR2_X1 U784 ( .A(n692), .B(n691), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n1002), .A2(G117), .ZN(n694) );
  NAND2_X1 U786 ( .A1(G129), .A2(n1003), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n1006), .A2(G141), .ZN(n695) );
  XOR2_X1 U789 ( .A(KEYINPUT94), .B(n695), .Z(n696) );
  NOR2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n993) );
  AND2_X1 U792 ( .A1(n993), .A2(G1996), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n924) );
  XNOR2_X1 U794 ( .A(KEYINPUT95), .B(n822), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n924), .A2(n702), .ZN(n813) );
  INV_X1 U796 ( .A(n813), .ZN(n713) );
  NAND2_X1 U797 ( .A1(G140), .A2(n1006), .ZN(n704) );
  NAND2_X1 U798 ( .A1(G104), .A2(n521), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U800 ( .A(KEYINPUT34), .B(n705), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n1002), .A2(G116), .ZN(n707) );
  NAND2_X1 U802 ( .A1(G128), .A2(n1003), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U804 ( .A(KEYINPUT35), .B(n708), .ZN(n709) );
  XNOR2_X1 U805 ( .A(KEYINPUT91), .B(n709), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U807 ( .A(KEYINPUT36), .B(n712), .ZN(n999) );
  XNOR2_X1 U808 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U809 ( .A1(n999), .A2(n819), .ZN(n926) );
  NAND2_X1 U810 ( .A1(n822), .A2(n926), .ZN(n817) );
  NAND2_X1 U811 ( .A1(n713), .A2(n817), .ZN(n808) );
  INV_X1 U812 ( .A(n841), .ZN(n1020) );
  INV_X1 U813 ( .A(n714), .ZN(n716) );
  INV_X1 U814 ( .A(n754), .ZN(n717) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n717), .ZN(n718) );
  XNOR2_X1 U816 ( .A(n718), .B(KEYINPUT26), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n754), .A2(G1341), .ZN(n720) );
  INV_X1 U818 ( .A(KEYINPUT100), .ZN(n719) );
  XNOR2_X1 U819 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U820 ( .A1(n1023), .A2(n721), .ZN(n722) );
  NAND2_X1 U821 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U822 ( .A(KEYINPUT64), .B(n724), .ZN(n730) );
  OR2_X1 U823 ( .A1(n1020), .A2(n730), .ZN(n729) );
  NAND2_X1 U824 ( .A1(G1348), .A2(n766), .ZN(n726) );
  NAND2_X1 U825 ( .A1(G2067), .A2(n717), .ZN(n725) );
  NAND2_X1 U826 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U827 ( .A(KEYINPUT101), .B(n727), .Z(n728) );
  NAND2_X1 U828 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U829 ( .A1(n1020), .A2(n730), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n741) );
  INV_X1 U831 ( .A(G2072), .ZN(n944) );
  NOR2_X1 U832 ( .A1(n754), .A2(n944), .ZN(n734) );
  XNOR2_X1 U833 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n733) );
  NAND2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n736) );
  OR2_X1 U835 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U836 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n766), .A2(G1956), .ZN(n737) );
  NAND2_X1 U838 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U839 ( .A(n739), .B(KEYINPUT99), .ZN(n742) );
  NAND2_X1 U840 ( .A1(n743), .A2(n742), .ZN(n740) );
  NAND2_X1 U841 ( .A1(n741), .A2(n740), .ZN(n746) );
  NOR2_X1 U842 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U843 ( .A(n744), .B(KEYINPUT28), .Z(n745) );
  NAND2_X1 U844 ( .A1(n746), .A2(n745), .ZN(n748) );
  XOR2_X1 U845 ( .A(G2078), .B(KEYINPUT25), .Z(n869) );
  NOR2_X1 U846 ( .A1(n869), .A2(n766), .ZN(n749) );
  XNOR2_X1 U847 ( .A(n749), .B(KEYINPUT97), .ZN(n751) );
  OR2_X1 U848 ( .A1(G1961), .A2(n717), .ZN(n750) );
  NAND2_X1 U849 ( .A1(n751), .A2(n750), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n760), .A2(G171), .ZN(n752) );
  NAND2_X1 U851 ( .A1(n753), .A2(n752), .ZN(n765) );
  NAND2_X1 U852 ( .A1(G8), .A2(n766), .ZN(n802) );
  NOR2_X1 U853 ( .A1(G1966), .A2(n802), .ZN(n779) );
  INV_X1 U854 ( .A(KEYINPUT96), .ZN(n756) );
  NOR2_X1 U855 ( .A1(G2084), .A2(n754), .ZN(n755) );
  XNOR2_X1 U856 ( .A(n756), .B(n755), .ZN(n775) );
  NAND2_X1 U857 ( .A1(G8), .A2(n775), .ZN(n757) );
  NOR2_X1 U858 ( .A1(n779), .A2(n757), .ZN(n758) );
  XOR2_X1 U859 ( .A(KEYINPUT30), .B(n758), .Z(n759) );
  NOR2_X1 U860 ( .A1(G168), .A2(n759), .ZN(n762) );
  NOR2_X1 U861 ( .A1(G171), .A2(n760), .ZN(n761) );
  XOR2_X1 U862 ( .A(KEYINPUT31), .B(n763), .Z(n764) );
  NAND2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n777), .A2(G286), .ZN(n771) );
  NOR2_X1 U865 ( .A1(G1971), .A2(n802), .ZN(n768) );
  NOR2_X1 U866 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U867 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U868 ( .A1(n769), .A2(G303), .ZN(n770) );
  NAND2_X1 U869 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U870 ( .A(n772), .B(KEYINPUT102), .ZN(n773) );
  NAND2_X1 U871 ( .A1(n773), .A2(G8), .ZN(n774) );
  XNOR2_X1 U872 ( .A(n774), .B(KEYINPUT32), .ZN(n783) );
  INV_X1 U873 ( .A(n775), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n776), .A2(G8), .ZN(n781) );
  INV_X1 U875 ( .A(n777), .ZN(n778) );
  NOR2_X1 U876 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n798) );
  NOR2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n850) );
  NOR2_X1 U880 ( .A1(G1971), .A2(G303), .ZN(n784) );
  NOR2_X1 U881 ( .A1(n850), .A2(n784), .ZN(n786) );
  INV_X1 U882 ( .A(KEYINPUT33), .ZN(n785) );
  AND2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n798), .A2(n787), .ZN(n791) );
  INV_X1 U885 ( .A(n802), .ZN(n788) );
  NAND2_X1 U886 ( .A1(G1976), .A2(G288), .ZN(n851) );
  AND2_X1 U887 ( .A1(n788), .A2(n851), .ZN(n789) );
  OR2_X1 U888 ( .A1(KEYINPUT33), .A2(n789), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U890 ( .A1(n850), .A2(KEYINPUT33), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n792), .A2(n802), .ZN(n793) );
  XOR2_X1 U892 ( .A(G1981), .B(G305), .Z(n838) );
  NAND2_X1 U893 ( .A1(n795), .A2(n838), .ZN(n806) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n796) );
  NAND2_X1 U895 ( .A1(G8), .A2(n796), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n799), .A2(n802), .ZN(n804) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U899 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  OR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  AND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  AND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n825) );
  XOR2_X1 U904 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n816) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n993), .ZN(n921) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U907 ( .A1(n866), .A2(n998), .ZN(n929) );
  NOR2_X1 U908 ( .A1(n811), .A2(n929), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n921), .A2(n814), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n816), .B(n815), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n819), .A2(n999), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n820), .B(KEYINPUT104), .ZN(n934) );
  NAND2_X1 U915 ( .A1(n821), .A2(n934), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U925 ( .A(G171), .ZN(G301) );
  NAND2_X1 U926 ( .A1(G136), .A2(n1006), .ZN(n832) );
  NAND2_X1 U927 ( .A1(G112), .A2(n1002), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n837) );
  NAND2_X1 U929 ( .A1(G124), .A2(n1003), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n833), .B(KEYINPUT44), .ZN(n835) );
  NAND2_X1 U931 ( .A1(G100), .A2(n521), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n835), .A2(n834), .ZN(n836) );
  NOR2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G162) );
  XNOR2_X1 U934 ( .A(G16), .B(KEYINPUT56), .ZN(n862) );
  XNOR2_X1 U935 ( .A(G1966), .B(G168), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n840), .B(KEYINPUT57), .ZN(n846) );
  XNOR2_X1 U938 ( .A(G1348), .B(KEYINPUT117), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n844) );
  XNOR2_X1 U940 ( .A(G1961), .B(G301), .ZN(n843) );
  NOR2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n848) );
  XNOR2_X1 U943 ( .A(G1341), .B(n1023), .ZN(n847) );
  NOR2_X1 U944 ( .A1(n848), .A2(n847), .ZN(n860) );
  XNOR2_X1 U945 ( .A(G1971), .B(G166), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(KEYINPUT118), .ZN(n856) );
  INV_X1 U947 ( .A(n850), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n854) );
  XNOR2_X1 U949 ( .A(G1956), .B(G299), .ZN(n853) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U952 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U953 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U954 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U955 ( .A(n863), .B(KEYINPUT119), .ZN(n888) );
  XOR2_X1 U956 ( .A(G34), .B(KEYINPUT116), .Z(n865) );
  XNOR2_X1 U957 ( .A(G2084), .B(KEYINPUT54), .ZN(n864) );
  XNOR2_X1 U958 ( .A(n865), .B(n864), .ZN(n884) );
  XNOR2_X1 U959 ( .A(G2090), .B(G35), .ZN(n882) );
  XNOR2_X1 U960 ( .A(G25), .B(n866), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n867), .A2(G28), .ZN(n868) );
  XOR2_X1 U962 ( .A(KEYINPUT113), .B(n868), .Z(n879) );
  XNOR2_X1 U963 ( .A(G33), .B(n944), .ZN(n873) );
  XNOR2_X1 U964 ( .A(G2067), .B(G26), .ZN(n871) );
  XNOR2_X1 U965 ( .A(G27), .B(n869), .ZN(n870) );
  NOR2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U967 ( .A1(n873), .A2(n872), .ZN(n876) );
  XNOR2_X1 U968 ( .A(KEYINPUT114), .B(G1996), .ZN(n874) );
  XNOR2_X1 U969 ( .A(G32), .B(n874), .ZN(n875) );
  NOR2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U971 ( .A(n877), .B(KEYINPUT115), .ZN(n878) );
  NOR2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT53), .B(n880), .ZN(n881) );
  NOR2_X1 U974 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U975 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U976 ( .A(KEYINPUT55), .B(n885), .ZN(n886) );
  NOR2_X1 U977 ( .A1(n886), .A2(G29), .ZN(n887) );
  NOR2_X1 U978 ( .A1(n888), .A2(n887), .ZN(n889) );
  NAND2_X1 U979 ( .A1(G11), .A2(n889), .ZN(n918) );
  XNOR2_X1 U980 ( .A(G20), .B(G1956), .ZN(n890) );
  XNOR2_X1 U981 ( .A(n890), .B(KEYINPUT121), .ZN(n896) );
  XNOR2_X1 U982 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n891) );
  XNOR2_X1 U983 ( .A(n891), .B(G4), .ZN(n892) );
  XNOR2_X1 U984 ( .A(G1348), .B(n892), .ZN(n894) );
  XNOR2_X1 U985 ( .A(G1981), .B(G6), .ZN(n893) );
  NOR2_X1 U986 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U987 ( .A1(n896), .A2(n895), .ZN(n899) );
  XNOR2_X1 U988 ( .A(KEYINPUT122), .B(G1341), .ZN(n897) );
  XNOR2_X1 U989 ( .A(G19), .B(n897), .ZN(n898) );
  NOR2_X1 U990 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U991 ( .A(KEYINPUT124), .B(n900), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n901), .B(KEYINPUT60), .ZN(n905) );
  XNOR2_X1 U993 ( .A(G1966), .B(G21), .ZN(n903) );
  XNOR2_X1 U994 ( .A(G1961), .B(G5), .ZN(n902) );
  NOR2_X1 U995 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U996 ( .A1(n905), .A2(n904), .ZN(n912) );
  XNOR2_X1 U997 ( .A(G1986), .B(G24), .ZN(n907) );
  XNOR2_X1 U998 ( .A(G1971), .B(G22), .ZN(n906) );
  NOR2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n909) );
  XOR2_X1 U1000 ( .A(G1976), .B(G23), .Z(n908) );
  NAND2_X1 U1001 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(KEYINPUT58), .B(n910), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1004 ( .A(KEYINPUT61), .B(n913), .Z(n915) );
  XNOR2_X1 U1005 ( .A(KEYINPUT120), .B(G16), .ZN(n914) );
  NOR2_X1 U1006 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1007 ( .A(KEYINPUT125), .B(n916), .Z(n917) );
  NOR2_X1 U1008 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1009 ( .A(n919), .B(KEYINPUT126), .ZN(n956) );
  XOR2_X1 U1010 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1011 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1012 ( .A(KEYINPUT51), .B(n922), .Z(n923) );
  NAND2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n932) );
  XOR2_X1 U1014 ( .A(G160), .B(G2084), .Z(n925) );
  NOR2_X1 U1015 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1016 ( .A1(n927), .A2(n1013), .ZN(n928) );
  NOR2_X1 U1017 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1018 ( .A(KEYINPUT111), .B(n930), .ZN(n931) );
  NOR2_X1 U1019 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1020 ( .A1(n934), .A2(n933), .ZN(n950) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n946) );
  NAND2_X1 U1022 ( .A1(n1006), .A2(G139), .ZN(n935) );
  XOR2_X1 U1023 ( .A(KEYINPUT107), .B(n935), .Z(n937) );
  NAND2_X1 U1024 ( .A1(n521), .A2(G103), .ZN(n936) );
  NAND2_X1 U1025 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1026 ( .A(KEYINPUT108), .B(n938), .ZN(n943) );
  NAND2_X1 U1027 ( .A1(n1002), .A2(G115), .ZN(n940) );
  NAND2_X1 U1028 ( .A1(G127), .A2(n1003), .ZN(n939) );
  NAND2_X1 U1029 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1030 ( .A(KEYINPUT47), .B(n941), .Z(n942) );
  NOR2_X1 U1031 ( .A1(n943), .A2(n942), .ZN(n994) );
  XNOR2_X1 U1032 ( .A(n944), .B(n994), .ZN(n945) );
  NOR2_X1 U1033 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1034 ( .A(KEYINPUT50), .B(n947), .Z(n948) );
  XNOR2_X1 U1035 ( .A(KEYINPUT112), .B(n948), .ZN(n949) );
  NOR2_X1 U1036 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n951), .ZN(n953) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n952) );
  NAND2_X1 U1039 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1040 ( .A1(n954), .A2(G29), .ZN(n955) );
  NAND2_X1 U1041 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1042 ( .A(KEYINPUT62), .B(n957), .Z(G311) );
  XNOR2_X1 U1043 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NOR2_X1 U1044 ( .A1(G860), .A2(n958), .ZN(n959) );
  XOR2_X1 U1045 ( .A(n960), .B(n959), .Z(G145) );
  INV_X1 U1046 ( .A(G120), .ZN(G236) );
  INV_X1 U1047 ( .A(G96), .ZN(G221) );
  INV_X1 U1048 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1049 ( .A1(n962), .A2(n961), .ZN(G325) );
  INV_X1 U1050 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1051 ( .A(G1976), .B(G2474), .ZN(n972) );
  XOR2_X1 U1052 ( .A(G1981), .B(G1966), .Z(n964) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G1986), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(n964), .B(n963), .ZN(n968) );
  XOR2_X1 U1055 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n966) );
  XNOR2_X1 U1056 ( .A(G1991), .B(G1956), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1058 ( .A(n968), .B(n967), .Z(n970) );
  XNOR2_X1 U1059 ( .A(G1961), .B(G1971), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n970), .B(n969), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n972), .B(n971), .ZN(G229) );
  XOR2_X1 U1062 ( .A(G2100), .B(G2096), .Z(n974) );
  XNOR2_X1 U1063 ( .A(G2072), .B(G2090), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n974), .B(n973), .ZN(n978) );
  XOR2_X1 U1065 ( .A(G2678), .B(KEYINPUT42), .Z(n976) );
  XNOR2_X1 U1066 ( .A(G2067), .B(KEYINPUT43), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1068 ( .A(n978), .B(n977), .Z(n980) );
  XNOR2_X1 U1069 ( .A(G2078), .B(G2084), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n980), .B(n979), .ZN(G227) );
  XNOR2_X1 U1071 ( .A(G1348), .B(G2454), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n981), .B(G2430), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n982), .B(G1341), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G2443), .B(G2427), .Z(n984) );
  XNOR2_X1 U1075 ( .A(G2438), .B(G2446), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n984), .B(n983), .ZN(n986) );
  XOR2_X1 U1077 ( .A(G2451), .B(G2435), .Z(n985) );
  XNOR2_X1 U1078 ( .A(n986), .B(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n988), .B(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n989), .A2(G14), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT105), .B(n990), .ZN(G401) );
  XOR2_X1 U1082 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n992) );
  XNOR2_X1 U1083 ( .A(G160), .B(KEYINPUT109), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n992), .B(n991), .ZN(n997) );
  XOR2_X1 U1085 ( .A(G164), .B(n993), .Z(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n997), .B(n996), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n999), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1001), .B(n1000), .ZN(n1017) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(G118), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(G130), .A2(n1003), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  NAND2_X1 U1093 ( .A1(G142), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1094 ( .A1(G106), .A2(n521), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(n1010), .B(KEYINPUT45), .Z(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(G162), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1100 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NOR2_X1 U1101 ( .A1(G37), .A2(n1018), .ZN(G395) );
  XOR2_X1 U1102 ( .A(n1019), .B(G286), .Z(n1022) );
  XNOR2_X1 U1103 ( .A(G171), .B(n1020), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(n1022), .B(n1021), .ZN(n1024) );
  XOR2_X1 U1105 ( .A(n1024), .B(n1023), .Z(n1025) );
  NOR2_X1 U1106 ( .A1(G37), .A2(n1025), .ZN(G397) );
  XNOR2_X1 U1107 ( .A(KEYINPUT110), .B(KEYINPUT49), .ZN(n1027) );
  NOR2_X1 U1108 ( .A1(G229), .A2(G227), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(n1027), .B(n1026), .ZN(n1029) );
  OR2_X1 U1110 ( .A1(n1032), .A2(G401), .ZN(n1028) );
  NOR2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  NOR2_X1 U1112 ( .A1(G395), .A2(G397), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(G225) );
  INV_X1 U1114 ( .A(G225), .ZN(G308) );
  INV_X1 U1115 ( .A(n1032), .ZN(G319) );
  INV_X1 U1116 ( .A(G108), .ZN(G238) );
endmodule

