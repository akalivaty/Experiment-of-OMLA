//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT78), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G107), .ZN(new_n193));
  OAI21_X1  g007(.A(G101), .B1(new_n193), .B2(KEYINPUT78), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(G104), .B2(new_n190), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n191), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n190), .A3(G104), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n203), .A2(new_n201), .A3(new_n200), .A4(new_n193), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT2), .B(G113), .Z(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n210), .A2(KEYINPUT5), .A3(G119), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(KEYINPUT80), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(KEYINPUT80), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(G113), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n209), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n198), .A2(new_n201), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT4), .B1(new_n217), .B2(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(new_n205), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(G101), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(KEYINPUT4), .ZN(new_n222));
  XOR2_X1   g036(.A(G116), .B(G119), .Z(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT2), .B(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n225), .A2(new_n209), .A3(KEYINPUT68), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n225), .B2(new_n209), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n216), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G110), .B(G122), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n216), .B(new_n231), .C1(new_n222), .C2(new_n229), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT6), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G143), .ZN(new_n238));
  INV_X1    g052(.A(G143), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT66), .B1(new_n239), .B2(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(G146), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g057(.A(G128), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n237), .A2(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(G146), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n243), .A4(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G125), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT0), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(KEYINPUT0), .B2(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n239), .A2(KEYINPUT66), .A3(G146), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n236), .B1(new_n237), .B2(G143), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n246), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n246), .A2(new_n247), .ZN(new_n265));
  OAI22_X1  g079(.A1(new_n261), .A2(new_n264), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n251), .B1(new_n250), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G224), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI221_X1 g084(.A(new_n251), .B1(new_n268), .B2(G953), .C1(new_n250), .C2(new_n266), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n230), .A2(new_n273), .A3(new_n232), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n235), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  OR3_X1    g091(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n269), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n231), .B(KEYINPUT8), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n206), .A2(new_n209), .A3(new_n215), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n206), .B1(new_n209), .B2(new_n215), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n283), .B2(new_n234), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n187), .B1(new_n275), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n275), .A2(new_n284), .A3(new_n187), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT79), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(KEYINPUT81), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n275), .A2(new_n284), .A3(new_n187), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(new_n285), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n295), .B2(new_n290), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(G234), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT22), .B(G137), .Z(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT75), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT70), .B(G953), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G221), .ZN(new_n305));
  INV_X1    g119(.A(G234), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n302), .B(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n310));
  INV_X1    g124(.A(G119), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(G128), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n312), .B(new_n313), .C1(G119), .C2(new_n253), .ZN(new_n314));
  XNOR2_X1  g128(.A(G119), .B(G128), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT24), .B(G110), .Z(new_n316));
  AOI22_X1  g130(.A1(new_n314), .A2(G110), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n250), .A2(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n250), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  AOI21_X1  g136(.A(G146), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n323), .A2(KEYINPUT72), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n322), .A3(G146), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n323), .B2(KEYINPUT72), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n317), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n314), .A2(G110), .B1(new_n315), .B2(new_n316), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n320), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n331), .B2(new_n237), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n330), .A2(KEYINPUT73), .A3(G146), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n328), .B(new_n325), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n327), .A2(KEYINPUT74), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT74), .B1(new_n327), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n309), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n327), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n308), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT25), .B1(new_n340), .B2(new_n299), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n342), .B(G902), .C1(new_n337), .C2(new_n339), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n300), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n300), .A2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n303), .A2(G210), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT27), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G101), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT69), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n226), .B2(new_n227), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n225), .A2(new_n209), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n225), .A2(new_n209), .A3(KEYINPUT68), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT69), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT11), .ZN(new_n362));
  INV_X1    g176(.A(G134), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(G137), .ZN(new_n364));
  INV_X1    g178(.A(G137), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT11), .A3(G134), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(G137), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G131), .ZN(new_n369));
  INV_X1    g183(.A(G131), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n364), .A2(new_n366), .A3(new_n370), .A4(new_n367), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n265), .A2(new_n258), .ZN(new_n375));
  INV_X1    g189(.A(new_n261), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n242), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n365), .A2(G134), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n370), .B1(new_n381), .B2(new_n367), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n245), .B2(new_n248), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n374), .A2(new_n377), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n361), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT28), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n361), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n228), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n353), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n361), .A2(new_n384), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n380), .A2(new_n383), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n266), .B1(new_n380), .B2(new_n369), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT30), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n384), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n393), .B1(new_n399), .B2(new_n228), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT31), .A3(new_n353), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n374), .A2(new_n377), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n380), .A2(new_n383), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n402), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n397), .B1(new_n402), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n228), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n385), .A3(new_n353), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT31), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n392), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(G472), .A2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n348), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n389), .A2(new_n391), .ZN(new_n414));
  INV_X1    g228(.A(new_n353), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT31), .B1(new_n400), .B2(new_n353), .ZN(new_n417));
  AND4_X1   g231(.A1(KEYINPUT31), .A2(new_n406), .A3(new_n385), .A4(new_n353), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT71), .A3(new_n411), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT32), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G472), .ZN(new_n423));
  INV_X1    g237(.A(new_n388), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n387), .B1(new_n361), .B2(new_n384), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n391), .B(new_n353), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT29), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(new_n353), .C2(new_n400), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n361), .A2(new_n384), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n386), .B2(new_n388), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n415), .A2(new_n427), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n423), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n401), .A2(new_n409), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n412), .B1(new_n434), .B2(new_n416), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(KEYINPUT32), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n347), .B1(new_n422), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G952), .ZN(new_n438));
  AOI211_X1 g252(.A(G953), .B(new_n438), .C1(G234), .C2(G237), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n304), .B(G902), .C1(new_n306), .C2(new_n349), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT87), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(G898), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n239), .A2(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n253), .A2(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G134), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n449), .A3(new_n363), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G116), .B(G122), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G122), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G116), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n190), .B1(new_n458), .B2(KEYINPUT14), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n190), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n453), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n239), .A2(KEYINPUT13), .A3(G128), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT83), .A3(new_n449), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT13), .B1(new_n239), .B2(G128), .ZN(new_n465));
  OAI221_X1 g279(.A(G134), .B1(KEYINPUT83), .B2(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n448), .A2(new_n449), .A3(new_n363), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n210), .A2(G122), .ZN(new_n468));
  OAI21_X1  g282(.A(G107), .B1(new_n458), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n462), .A2(KEYINPUT84), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n453), .A2(new_n460), .A3(new_n472), .A4(new_n461), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT9), .B(G234), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n474), .A2(new_n298), .A3(G953), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n363), .B1(new_n448), .B2(new_n449), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n461), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n210), .A2(G122), .ZN(new_n479));
  OAI21_X1  g293(.A(G107), .B1(new_n479), .B2(new_n455), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n455), .B2(new_n454), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT84), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n466), .A2(new_n470), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n473), .ZN(new_n484));
  INV_X1    g298(.A(new_n475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n476), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n447), .B1(new_n487), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n476), .A2(new_n486), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT85), .A3(new_n299), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n446), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT85), .B1(new_n489), .B2(new_n299), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n445), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT86), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n447), .B(G902), .C1(new_n476), .C2(new_n486), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n445), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n488), .A2(new_n446), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n443), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n303), .A2(G143), .A3(G214), .A4(new_n349), .ZN(new_n502));
  OR2_X1    g316(.A1(KEYINPUT70), .A2(G953), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT70), .A2(G953), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n503), .A2(G214), .A3(new_n349), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n239), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n370), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(new_n370), .A3(new_n506), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n502), .A2(new_n506), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT17), .A3(G131), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n324), .A2(new_n326), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n516), .A3(KEYINPUT17), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n511), .A2(new_n514), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G113), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n188), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(KEYINPUT18), .A3(G131), .ZN(new_n521));
  OAI22_X1  g335(.A1(new_n332), .A2(new_n333), .B1(new_n237), .B2(new_n331), .ZN(new_n522));
  NAND2_X1  g336(.A1(KEYINPUT18), .A2(G131), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n502), .A2(new_n506), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n520), .ZN(new_n527));
  INV_X1    g341(.A(new_n525), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n330), .B(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n325), .B1(new_n529), .B2(G146), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n508), .B2(new_n510), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G475), .A2(G902), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n501), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  AOI211_X1 g350(.A(KEYINPUT20), .B(new_n536), .C1(new_n526), .C2(new_n532), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n518), .A2(new_n525), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n527), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n539), .B2(new_n526), .ZN(new_n540));
  INV_X1    g354(.A(G475), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n535), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n500), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n474), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n305), .B1(new_n545), .B2(new_n299), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT4), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n219), .B2(new_n220), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n377), .B1(new_n549), .B2(new_n218), .ZN(new_n550));
  INV_X1    g364(.A(new_n374), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n244), .A2(new_n265), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n248), .ZN(new_n553));
  INV_X1    g367(.A(new_n195), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n245), .B2(new_n248), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n557), .A2(new_n558), .B1(new_n206), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n550), .A2(new_n551), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n557), .B1(new_n249), .B2(new_n206), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n562), .A2(KEYINPUT12), .A3(new_n374), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT12), .B1(new_n562), .B2(new_n374), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n303), .A2(G227), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT76), .ZN(new_n567));
  XNOR2_X1  g381(.A(G110), .B(G140), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n550), .A2(new_n560), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n374), .ZN(new_n572));
  INV_X1    g386(.A(new_n569), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n561), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(G469), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(G469), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n550), .A2(new_n551), .A3(new_n560), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n551), .B1(new_n550), .B2(new_n560), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n569), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n561), .B(new_n573), .C1(new_n563), .C2(new_n564), .ZN(new_n581));
  AOI211_X1 g395(.A(G469), .B(G902), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n547), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n544), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n297), .A2(new_n437), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  OAI21_X1  g400(.A(G472), .B1(new_n410), .B2(G902), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n413), .A2(new_n587), .A3(new_n420), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n588), .A2(new_n347), .A3(new_n583), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n444), .A2(new_n299), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n487), .A2(G902), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n444), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n489), .A2(KEYINPUT33), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n489), .A2(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(G478), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n542), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n443), .ZN(new_n599));
  INV_X1    g413(.A(new_n289), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n295), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n589), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  AND2_X1   g418(.A1(new_n526), .A2(new_n532), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT20), .B1(new_n605), .B2(new_n536), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT88), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n533), .A2(new_n501), .A3(new_n534), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT88), .B1(new_n535), .B2(new_n537), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n540), .A2(new_n541), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n494), .A2(new_n499), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n443), .B(KEYINPUT89), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n610), .A2(new_n611), .ZN(new_n618));
  INV_X1    g432(.A(new_n499), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n498), .B1(new_n496), .B2(new_n497), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n618), .A2(new_n621), .A3(new_n609), .A4(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT90), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n589), .A2(new_n601), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  OR2_X1    g440(.A1(new_n335), .A2(new_n336), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n309), .A2(KEYINPUT36), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n345), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n344), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n588), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n297), .A2(new_n584), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  AOI21_X1  g451(.A(new_n583), .B1(new_n422), .B2(new_n436), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n288), .A2(new_n289), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n633), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n439), .B1(new_n441), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n612), .A2(new_n613), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n638), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  NAND2_X1  g459(.A1(new_n621), .A2(new_n542), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n633), .A2(new_n289), .ZN(new_n647));
  INV_X1    g461(.A(new_n583), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT92), .B(KEYINPUT39), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n642), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n646), .B(new_n647), .C1(new_n651), .C2(KEYINPUT40), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n400), .A2(new_n415), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n393), .A2(new_n429), .A3(new_n353), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(G902), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n423), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n435), .B2(KEYINPUT32), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n422), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n295), .B(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n652), .A2(new_n658), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT93), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  INV_X1    g478(.A(KEYINPUT94), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n598), .B2(new_n642), .ZN(new_n666));
  INV_X1    g480(.A(new_n642), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n542), .A2(new_n597), .A3(KEYINPUT94), .A4(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n638), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  NAND2_X1  g485(.A1(new_n422), .A2(new_n436), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n580), .A2(new_n581), .ZN(new_n673));
  OAI21_X1  g487(.A(G469), .B1(new_n673), .B2(G902), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT95), .ZN(new_n675));
  INV_X1    g489(.A(new_n582), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(KEYINPUT95), .B(G469), .C1(new_n673), .C2(G902), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n546), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n347), .A2(new_n598), .A3(new_n443), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n672), .A2(new_n679), .A3(new_n601), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  INV_X1    g497(.A(new_n347), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n623), .A2(new_n617), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n672), .A2(new_n601), .A3(new_n679), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n210), .ZN(G18));
  AND3_X1   g502(.A1(new_n500), .A2(new_n543), .A3(new_n632), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n672), .A2(new_n679), .A3(new_n601), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  OAI22_X1  g505(.A1(new_n417), .A2(new_n418), .B1(new_n353), .B2(new_n430), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n411), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n684), .A2(new_n587), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n621), .A2(new_n542), .A3(new_n616), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n679), .A3(new_n601), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  NAND2_X1  g511(.A1(new_n666), .A2(new_n668), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n587), .A2(new_n693), .A3(new_n632), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT96), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n587), .A2(new_n693), .A3(new_n632), .A4(KEYINPUT96), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n679), .A2(new_n601), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  INV_X1    g520(.A(KEYINPUT97), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n583), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n294), .A2(new_n285), .A3(new_n600), .ZN(new_n709));
  OAI211_X1 g523(.A(KEYINPUT97), .B(new_n547), .C1(new_n577), .C2(new_n582), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT98), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n708), .A2(new_n709), .A3(new_n713), .A4(new_n710), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n421), .B1(new_n410), .B2(new_n412), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n347), .B1(new_n436), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n717), .A3(KEYINPUT42), .A4(new_n669), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT99), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n715), .A2(new_n720), .A3(new_n437), .A4(new_n669), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n672), .A2(new_n684), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n714), .B2(new_n712), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n720), .B1(new_n725), .B2(new_n669), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT100), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n715), .A2(new_n437), .A3(new_n669), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT100), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n722), .A4(new_n721), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n719), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n370), .ZN(G33));
  NAND2_X1  g547(.A1(new_n725), .A2(new_n643), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT102), .B(G134), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G36));
  AND2_X1   g552(.A1(new_n570), .A2(new_n574), .ZN(new_n739));
  OAI21_X1  g553(.A(G469), .B1(new_n739), .B2(KEYINPUT45), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n576), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n676), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(KEYINPUT105), .B(new_n676), .C1(new_n746), .C2(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n746), .A2(new_n747), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n547), .A3(new_n650), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n542), .A2(new_n596), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT43), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n588), .A3(new_n632), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT107), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  INV_X1    g576(.A(new_n709), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n762), .A2(KEYINPUT106), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT106), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT108), .B(G137), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G39));
  NOR4_X1   g583(.A1(new_n672), .A2(new_n698), .A3(new_n684), .A4(new_n763), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n753), .A2(KEYINPUT47), .A3(new_n547), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT47), .B1(new_n753), .B2(new_n547), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n776), .B(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT110), .B(G140), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G42));
  NAND3_X1  g594(.A1(new_n757), .A2(new_n694), .A3(new_n439), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n661), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n600), .A3(new_n783), .A4(new_n679), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT50), .Z(new_n785));
  AND3_X1   g599(.A1(new_n679), .A2(new_n439), .A3(new_n709), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n757), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n701), .B2(new_n702), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n658), .A2(new_n347), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n542), .A2(new_n597), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n785), .A2(new_n792), .A3(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n753), .A2(new_n547), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n677), .A2(new_n678), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n546), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n771), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT117), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n781), .A2(new_n763), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n799), .A2(KEYINPUT117), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n793), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n786), .A2(new_n717), .A3(new_n757), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n790), .A2(new_n542), .A3(new_n597), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n438), .B(G953), .C1(new_n782), .C2(new_n704), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n785), .A2(new_n792), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n772), .B2(new_n773), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n796), .A2(KEYINPUT116), .A3(new_n771), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n798), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n811), .B1(new_n815), .B2(new_n801), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n804), .B(new_n810), .C1(new_n816), .C2(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n727), .A2(new_n731), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n718), .ZN(new_n819));
  INV_X1    g633(.A(new_n736), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n715), .A2(new_n703), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n632), .A2(new_n496), .A3(new_n497), .A4(new_n667), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n612), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n638), .A2(new_n709), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n542), .B1(new_n496), .B2(new_n497), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(KEYINPUT112), .B2(new_n598), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(KEYINPUT112), .B2(new_n598), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n297), .A3(new_n589), .A4(new_n616), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n585), .A3(new_n635), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n681), .A2(new_n696), .A3(new_n690), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n687), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT111), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n831), .B2(new_n687), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n825), .B(new_n830), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n638), .B(new_n640), .C1(new_n669), .C2(new_n643), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n633), .A2(new_n667), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n839), .B2(new_n583), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n639), .A2(new_n646), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n648), .A2(KEYINPUT113), .A3(new_n633), .A4(new_n667), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n658), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n705), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n705), .A2(KEYINPUT52), .A3(new_n837), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n819), .A2(new_n820), .A3(new_n836), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g663(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n850));
  AOI21_X1  g664(.A(new_n736), .B1(new_n818), .B2(new_n718), .ZN(new_n851));
  INV_X1    g665(.A(new_n830), .ZN(new_n852));
  INV_X1    g666(.A(new_n825), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT53), .A4(new_n832), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n844), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n844), .A2(new_n855), .A3(KEYINPUT52), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n831), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n685), .A2(new_n686), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT111), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n831), .A2(new_n687), .A3(new_n834), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n853), .B(new_n852), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n732), .A2(new_n736), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n857), .A2(new_n858), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n846), .A2(new_n847), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n732), .A2(new_n867), .A3(new_n736), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n850), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n862), .B1(new_n874), .B2(new_n861), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n817), .A2(new_n875), .B1(G952), .B2(G953), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n797), .B(KEYINPUT49), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n542), .A2(new_n596), .A3(new_n290), .A4(new_n546), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n783), .A3(new_n789), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n303), .A2(G952), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n860), .A2(new_n299), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(G210), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n235), .A2(new_n274), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT119), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n272), .B(KEYINPUT55), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(KEYINPUT120), .A3(KEYINPUT121), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n885), .B(new_n886), .C1(new_n883), .C2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n881), .B1(new_n892), .B2(new_n894), .ZN(G51));
  NAND2_X1  g709(.A1(new_n851), .A2(new_n859), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n872), .B2(new_n873), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(G902), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n745), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n860), .B2(new_n861), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(KEYINPUT122), .A3(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n862), .A3(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n576), .B(KEYINPUT57), .Z(new_n904));
  AOI21_X1  g718(.A(new_n673), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n905), .B2(KEYINPUT123), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n907));
  INV_X1    g721(.A(new_n904), .ZN(new_n908));
  AOI221_X4 g722(.A(KEYINPUT54), .B1(new_n851), .B2(new_n859), .C1(new_n849), .C2(new_n850), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n911), .B2(new_n902), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n912), .B2(new_n673), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n881), .B1(new_n906), .B2(new_n913), .ZN(G54));
  NAND4_X1  g728(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .A4(new_n533), .ZN(new_n915));
  NAND2_X1  g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n605), .B1(new_n898), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n881), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT124), .Z(G60));
  NAND2_X1  g734(.A1(new_n593), .A2(new_n594), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n590), .B(KEYINPUT59), .Z(new_n922));
  AND3_X1   g736(.A1(new_n903), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n875), .B2(new_n922), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n881), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT60), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n897), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n340), .B(KEYINPUT125), .Z(new_n929));
  AOI21_X1  g743(.A(new_n881), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n629), .A2(new_n630), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n928), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT126), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(KEYINPUT126), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT127), .Z(new_n936));
  AND3_X1   g750(.A1(new_n932), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n932), .B2(new_n934), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  OAI21_X1  g753(.A(G953), .B1(new_n442), .B2(new_n268), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n830), .B1(new_n833), .B2(new_n835), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n304), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n888), .B1(G898), .B2(new_n303), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  AND2_X1   g758(.A1(new_n841), .A2(new_n717), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n755), .B1(new_n766), .B2(new_n945), .ZN(new_n946));
  AND4_X1   g760(.A1(new_n705), .A2(new_n946), .A3(new_n851), .A4(new_n837), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n778), .A3(new_n303), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n399), .B(new_n529), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(G900), .B2(new_n304), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n663), .A2(new_n705), .A3(new_n837), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n651), .A2(new_n763), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n828), .A2(new_n437), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n767), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n775), .B2(new_n777), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n949), .B1(new_n957), .B2(new_n304), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n303), .B1(G227), .B2(G900), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n951), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n957), .B2(new_n941), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n918), .B1(new_n968), .B2(new_n653), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n400), .A2(new_n353), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n967), .B(new_n874), .C1(new_n407), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n400), .A2(new_n415), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n947), .A2(new_n778), .A3(new_n941), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n966), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n969), .A2(new_n971), .A3(new_n974), .ZN(G57));
endmodule


