//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n461), .B2(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n469), .B2(new_n462), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n470), .B2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n461), .A2(new_n462), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NOR2_X1   g062(.A1(new_n462), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n480), .A2(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n471), .A2(new_n472), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n462), .A3(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n498), .A2(KEYINPUT4), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n461), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n496), .B(new_n497), .C1(new_n501), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT6), .B1(KEYINPUT70), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  AND3_X1   g089(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n515), .A2(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OAI221_X1 g098(.A(new_n513), .B1(new_n514), .B2(new_n518), .C1(new_n519), .C2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  INV_X1    g100(.A(new_n518), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT71), .B(G51), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n512), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n516), .A2(new_n517), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n526), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n512), .A2(G52), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR3_X1    g121(.A1(new_n546), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n526), .A2(G81), .B1(new_n512), .B2(G43), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT72), .B1(new_n546), .B2(new_n519), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n510), .A2(new_n511), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n512), .A2(new_n561), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n538), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G651), .A2(new_n566), .B1(new_n526), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  OAI21_X1  g143(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n569));
  OAI211_X1 g144(.A(G49), .B(G543), .C1(new_n515), .C2(new_n509), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n518), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n557), .A2(KEYINPUT73), .A3(G87), .A4(new_n522), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  INV_X1    g154(.A(G73), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n538), .A2(new_n579), .B1(new_n580), .B2(new_n508), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n581), .B2(G651), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n512), .A2(G48), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n557), .A2(G86), .A3(new_n522), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n579), .B1(new_n520), .B2(new_n521), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n580), .A2(new_n508), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n578), .B(G651), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n583), .A2(new_n586), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n526), .A2(G85), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT75), .B(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n558), .B2(new_n592), .C1(new_n519), .C2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n518), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n538), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n512), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n596), .B1(new_n606), .B2(new_n595), .ZN(G284));
  AOI21_X1  g182(.A(new_n596), .B1(new_n606), .B2(new_n595), .ZN(G321));
  NOR2_X1   g183(.A1(G286), .A2(new_n595), .ZN(new_n609));
  XNOR2_X1  g184(.A(G299), .B(KEYINPUT77), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n595), .ZN(G297));
  AOI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(new_n595), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NOR2_X1   g189(.A1(new_n551), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n606), .A2(new_n613), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT78), .Z(G323));
  XOR2_X1   g193(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n619));
  XNOR2_X1  g194(.A(G323), .B(new_n619), .ZN(G282));
  NAND2_X1  g195(.A1(new_n461), .A2(new_n464), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(new_n626));
  OR3_X1    g201(.A1(new_n462), .A2(KEYINPUT82), .A3(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT82), .B1(new_n462), .B2(G111), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  AND4_X1   g204(.A1(G2104), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n480), .A2(G123), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT81), .Z(new_n632));
  NOR2_X1   g207(.A1(new_n498), .A2(G2105), .ZN(new_n633));
  AOI211_X1 g208(.A(new_n630), .B(new_n632), .C1(G135), .C2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n634), .A2(new_n635), .B1(new_n624), .B2(new_n623), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n626), .B(new_n636), .C1(new_n635), .C2(new_n634), .ZN(G156));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT84), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT83), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n643), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n643), .B(new_n650), .ZN(new_n654));
  INV_X1    g229(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n653), .A2(G14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g233(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n663), .B2(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n672), .A2(new_n673), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n686), .B(new_n685), .S(new_n679), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT90), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n684), .A2(new_n690), .A3(new_n687), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n689), .A2(new_n691), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n689), .B2(new_n691), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n551), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n700), .B2(G19), .ZN(new_n702));
  INV_X1    g277(.A(G1341), .ZN(new_n703));
  INV_X1    g278(.A(G2084), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(KEYINPUT24), .B2(G34), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(KEYINPUT24), .B2(G34), .ZN(new_n707));
  INV_X1    g282(.A(G160), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G29), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n702), .A2(new_n703), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(G32), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G129), .B2(new_n480), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n633), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(new_n705), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT27), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1996), .ZN(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G35), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G162), .B2(G29), .ZN(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT100), .B(KEYINPUT29), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n705), .A2(G27), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT99), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n705), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2078), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  NAND2_X1  g306(.A1(G171), .A2(G16), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT97), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n730), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n710), .A2(new_n720), .A3(new_n726), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n705), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n480), .A2(G128), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G116), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n633), .B2(G140), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(G29), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(G115), .A2(G2104), .ZN(new_n751));
  INV_X1    g326(.A(G127), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n498), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G2105), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n757), .C1(new_n758), .C2(new_n485), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n762));
  OAI21_X1  g337(.A(G29), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G33), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(G29), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n750), .B1(G2072), .B2(new_n765), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n766), .B1(new_n703), .B2(new_n702), .C1(G2072), .C2(new_n765), .ZN(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(KEYINPUT30), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT96), .ZN(new_n770));
  AOI211_X1 g345(.A(G29), .B(new_n770), .C1(KEYINPUT30), .C2(new_n768), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT31), .B(G11), .Z(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n634), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(new_n735), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n700), .A2(G21), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G286), .B2(G16), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n775), .A2(G1961), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n774), .B(new_n779), .C1(new_n776), .C2(new_n778), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n737), .B(new_n767), .C1(KEYINPUT98), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n700), .A2(G20), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT23), .Z(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT102), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT101), .B(G1956), .Z(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n709), .A2(new_n704), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  NOR4_X1   g367(.A1(new_n782), .A2(new_n789), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G4), .A2(G16), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n606), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n781), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT103), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n700), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n700), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(G6), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G305), .B2(new_n700), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  OAI21_X1  g382(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n576), .A2(new_n700), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n700), .B2(G23), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n810), .A2(new_n811), .B1(new_n806), .B2(new_n807), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n808), .A2(new_n813), .A3(KEYINPUT34), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT34), .B1(new_n808), .B2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n480), .A2(G119), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n462), .A2(G107), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n818));
  INV_X1    g393(.A(G131), .ZN(new_n819));
  OAI221_X1 g394(.A(new_n816), .B1(new_n817), .B2(new_n818), .C1(new_n819), .C2(new_n485), .ZN(new_n820));
  MUX2_X1   g395(.A(G25), .B(new_n820), .S(G29), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n700), .A2(G24), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G290), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT91), .B(G1986), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n814), .A2(new_n815), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n800), .A2(new_n835), .ZN(G150));
  INV_X1    g411(.A(G150), .ZN(G311));
  NAND2_X1  g412(.A1(new_n526), .A2(G93), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n512), .A2(G55), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n838), .B(new_n839), .C1(new_n519), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT104), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(KEYINPUT104), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n551), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n549), .A2(new_n550), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n606), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT105), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n841), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n747), .B(new_n716), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n633), .A2(G142), .B1(G130), .B2(new_n480), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n862));
  INV_X1    g437(.A(G118), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n861), .A2(new_n862), .B1(new_n863), .B2(G2105), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n862), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n859), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n761), .A2(KEYINPUT106), .A3(new_n762), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n760), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n506), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT106), .B1(new_n761), .B2(new_n762), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n870), .A3(new_n760), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(G164), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n820), .B(new_n622), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n873), .B2(new_n876), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n877), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n867), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G160), .B(G162), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n634), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n881), .A2(new_n885), .A3(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g468(.A(new_n848), .B(new_n616), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n604), .B(G299), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n604), .A2(G299), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n604), .A2(G299), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(KEYINPUT41), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n903), .B2(new_n894), .ZN(new_n904));
  XNOR2_X1  g479(.A(G305), .B(G290), .ZN(new_n905));
  XNOR2_X1  g480(.A(G303), .B(new_n576), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n904), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n841), .A2(new_n595), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  OAI21_X1  g491(.A(G286), .B1(G171), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(G301), .A2(KEYINPUT109), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n845), .A2(new_n846), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n845), .A2(new_n846), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n844), .A2(new_n847), .A3(new_n920), .A4(new_n919), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n903), .ZN(new_n927));
  INV_X1    g502(.A(new_n895), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G37), .B1(new_n930), .B2(new_n907), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  INV_X1    g507(.A(new_n907), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(new_n933), .A3(new_n929), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n902), .B1(new_n924), .B2(new_n925), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n907), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT44), .Z(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n501), .A2(new_n505), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n496), .A2(new_n497), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n466), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n462), .B1(new_n473), .B2(new_n467), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n475), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT67), .B(new_n462), .C1(new_n473), .C2(new_n467), .ZN(new_n953));
  OAI211_X1 g528(.A(G40), .B(new_n950), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT46), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT123), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n747), .A2(G2067), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n742), .A2(new_n749), .A3(new_n746), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n717), .B1(new_n963), .B2(G1996), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT124), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT47), .ZN(new_n968));
  INV_X1    g543(.A(new_n955), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n716), .B(new_n956), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n820), .A2(new_n823), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n820), .A2(new_n823), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n961), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n971), .A2(KEYINPUT48), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(KEYINPUT48), .B2(new_n971), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n961), .A2(new_n972), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n960), .B1(new_n978), .B2(new_n973), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n955), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT122), .Z(new_n981));
  NOR3_X1   g556(.A1(new_n968), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n466), .C1(new_n470), .C2(new_n476), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n490), .A2(new_n495), .B1(new_n480), .B2(G126), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT4), .B1(new_n498), .B2(new_n500), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n461), .A2(new_n502), .A3(new_n504), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(new_n985), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1956), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(G299), .A2(KEYINPUT57), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n563), .B2(new_n567), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n506), .B2(new_n944), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n954), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n948), .A2(G1384), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n506), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT56), .B(G2072), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n995), .A2(new_n999), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n954), .A2(new_n947), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n993), .A2(new_n796), .B1(new_n749), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n604), .B(KEYINPUT76), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n999), .B1(new_n995), .B2(new_n1005), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT114), .B(KEYINPUT61), .Z(new_n1013));
  AND3_X1   g588(.A1(new_n995), .A2(new_n999), .A3(new_n1005), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1007), .A2(new_n749), .ZN(new_n1016));
  AOI211_X1 g591(.A(KEYINPUT50), .B(G1384), .C1(new_n986), .C2(new_n989), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n991), .B1(new_n506), .B2(new_n944), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n954), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT60), .B(new_n1016), .C1(new_n1019), .C2(G1348), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n1009), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1008), .A2(new_n606), .A3(KEYINPUT60), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1019), .B2(G1348), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n995), .A2(new_n1005), .ZN(new_n1027));
  INV_X1    g602(.A(new_n999), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT61), .A3(new_n1006), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1015), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n949), .A2(new_n985), .A3(new_n956), .A4(new_n1003), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1001), .A2(KEYINPUT113), .A3(new_n956), .A4(new_n1003), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT58), .B(G1341), .Z(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n954), .B2(new_n947), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n551), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1012), .B1(new_n1031), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT115), .B(new_n1012), .C1(new_n1031), .C2(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2078), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G40), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n466), .A2(new_n951), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n949), .A2(new_n1003), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1019), .B2(G1961), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1002), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n986), .B2(new_n989), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1000), .A2(new_n954), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G2078), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G171), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n949), .A2(new_n985), .A3(new_n1058), .A4(new_n1003), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1049), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1003), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1056), .A2(KEYINPUT112), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n1001), .A3(new_n1050), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n993), .A2(new_n731), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1062), .A2(new_n1067), .A3(new_n1068), .A4(G301), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1060), .A2(KEYINPUT54), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n949), .A2(new_n985), .A3(new_n1003), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1019), .A2(new_n723), .B1(new_n1076), .B2(new_n803), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1981), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n583), .A2(new_n586), .A3(new_n1080), .A4(new_n589), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n589), .A2(new_n584), .A3(new_n585), .ZN(new_n1082));
  OAI21_X1  g657(.A(G1981), .B1(new_n1082), .B2(new_n582), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1083), .A3(KEYINPUT111), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n1085));
  NAND3_X1  g660(.A1(G305), .A2(new_n1085), .A3(G1981), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT49), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n954), .B2(new_n947), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1084), .A2(new_n1091), .A3(new_n1086), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT110), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n576), .A2(new_n1095), .A3(G1976), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n574), .A2(new_n575), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n569), .A2(new_n570), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G1976), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT110), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1094), .B1(new_n1101), .B2(new_n1090), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1094), .B1(new_n576), .B2(G1976), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1103), .A2(new_n1089), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n983), .A2(new_n985), .A3(new_n992), .A4(new_n723), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1057), .B2(G1971), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n1074), .A3(G8), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1079), .A2(new_n1093), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1070), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n1112));
  NAND3_X1  g687(.A1(new_n1062), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1062), .A2(new_n1068), .A3(G301), .A4(new_n1053), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(KEYINPUT119), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1118), .B(new_n1112), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1111), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G286), .A2(G8), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n949), .A2(new_n985), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1063), .B(new_n1055), .C1(new_n986), .C2(new_n989), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT112), .B1(new_n506), .B2(new_n1002), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n776), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1019), .A2(new_n704), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1078), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1121), .B1(new_n1129), .B2(KEYINPUT116), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1966), .B1(new_n1066), .B2(new_n1001), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n704), .A2(new_n983), .A3(new_n985), .A4(new_n992), .ZN(new_n1132));
  OAI21_X1  g707(.A(G8), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT51), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1121), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(KEYINPUT51), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1133), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1137), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1128), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1120), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1048), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G288), .A2(G1976), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1093), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1089), .B1(new_n1147), .B2(new_n1081), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1103), .A2(new_n1089), .A3(new_n1104), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT52), .B1(new_n1103), .B2(new_n1089), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1092), .A2(new_n1090), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1091), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(new_n1109), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1109), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1074), .B1(new_n1108), .B2(G8), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1153), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1133), .A2(G286), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1159), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1110), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1155), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT120), .B1(new_n1145), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1167), .B(new_n1164), .C1(new_n1048), .C2(new_n1144), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1143), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1128), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT51), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1138), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1129), .A2(KEYINPUT116), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1139), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT117), .B1(new_n1129), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1133), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1171), .B(new_n1173), .C1(new_n1177), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1169), .B1(new_n1172), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1173), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT62), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1186), .A2(KEYINPUT121), .A3(new_n1182), .A4(new_n1170), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1166), .A2(new_n1168), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(G290), .B(G1986), .Z(new_n1190));
  AOI21_X1  g765(.A(new_n969), .B1(new_n975), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n982), .B1(new_n1189), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(G319), .ZN(new_n1194));
  NOR3_X1   g768(.A1(new_n657), .A2(new_n1194), .A3(G227), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1195), .B1(new_n697), .B2(new_n698), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n890), .B2(new_n891), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n942), .A2(KEYINPUT126), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g772(.A(KEYINPUT126), .B1(new_n942), .B2(new_n1197), .ZN(new_n1199));
  NOR3_X1   g773(.A1(new_n1198), .A2(new_n1199), .A3(KEYINPUT127), .ZN(new_n1200));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n932), .B1(new_n931), .B2(new_n934), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n1203));
  OAI21_X1  g777(.A(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n942), .A2(KEYINPUT126), .A3(new_n1197), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1201), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n1200), .A2(new_n1208), .ZN(G308));
  NAND2_X1  g783(.A1(new_n1206), .A2(new_n1207), .ZN(G225));
endmodule


