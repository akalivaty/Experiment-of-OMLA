//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT74), .A3(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT3), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n194), .A2(new_n189), .A3(KEYINPUT74), .A4(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT4), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G101), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(KEYINPUT76), .A3(new_n197), .A4(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n204), .B(new_n206), .C1(new_n209), .C2(new_n210), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n196), .A2(G101), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT75), .B(G101), .Z(new_n216));
  NAND4_X1  g030(.A1(new_n216), .A2(new_n193), .A3(new_n191), .A4(new_n195), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT10), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n205), .B(G146), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n210), .A2(new_n203), .A3(G143), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n221), .A2(KEYINPUT65), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT65), .B1(new_n221), .B2(new_n222), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n204), .A3(new_n206), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n220), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n192), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n217), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n221), .A3(new_n222), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n228), .A2(new_n232), .B1(new_n220), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT11), .ZN(new_n236));
  INV_X1    g050(.A(G134), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(G137), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .A3(G134), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G131), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n241), .A3(new_n244), .A4(new_n239), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n219), .A2(new_n235), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n219), .A2(new_n235), .A3(KEYINPUT77), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G110), .B(G140), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n254), .A2(G227), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n253), .B(new_n255), .Z(new_n256));
  AOI21_X1  g070(.A(KEYINPUT78), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n258), .B(new_n259), .C1(new_n250), .C2(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n221), .A2(new_n222), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n221), .A2(KEYINPUT65), .A3(new_n222), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n227), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n234), .B1(new_n232), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n246), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n257), .A2(new_n260), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n247), .B1(new_n219), .B2(new_n235), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n256), .B1(new_n252), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n187), .B(new_n188), .C1(new_n269), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT79), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n252), .A2(new_n256), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n258), .ZN(new_n277));
  INV_X1    g091(.A(new_n268), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n252), .A2(KEYINPUT78), .A3(new_n256), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n272), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT79), .A3(new_n187), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n252), .A2(new_n256), .A3(new_n271), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n268), .B1(new_n250), .B2(new_n251), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n256), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n188), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n275), .A2(new_n283), .B1(G469), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G125), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n212), .B2(new_n213), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n289), .B2(new_n265), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT81), .B(G224), .Z(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n254), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n291), .B(new_n293), .Z(new_n294));
  XOR2_X1   g108(.A(G110), .B(G122), .Z(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(G116), .B(G119), .Z(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT2), .B(G113), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n202), .A2(new_n300), .A3(new_n218), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G116), .ZN(new_n305));
  OAI211_X1 g119(.A(G113), .B(new_n305), .C1(new_n297), .C2(new_n303), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n232), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n301), .A2(new_n307), .A3(new_n296), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(KEYINPUT6), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n309), .A2(new_n312), .A3(KEYINPUT6), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT6), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT80), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n294), .B(new_n311), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n291), .B1(new_n254), .B2(new_n292), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n317), .A2(KEYINPUT7), .B1(new_n291), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n306), .A2(new_n302), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n232), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n295), .B(KEYINPUT8), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n319), .B(new_n310), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n316), .A2(new_n188), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n325), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n316), .A2(new_n188), .A3(new_n329), .A4(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(G234), .A2(G237), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G952), .A3(new_n254), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT21), .B(G898), .Z(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(G902), .A3(G953), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G214), .B1(G237), .B2(G902), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n331), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT9), .B(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n188), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n341), .A2(G221), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(KEYINPUT16), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(KEYINPUT16), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n289), .A2(G140), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n346), .A3(KEYINPUT70), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n345), .A2(KEYINPUT70), .A3(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n352), .B2(KEYINPUT16), .ZN(new_n353));
  OAI211_X1 g167(.A(G146), .B(new_n347), .C1(new_n353), .C2(new_n344), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n350), .B2(new_n351), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT71), .B1(new_n357), .B2(new_n348), .ZN(new_n358));
  AOI21_X1  g172(.A(G146), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n343), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n347), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n203), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT87), .A3(new_n354), .ZN(new_n363));
  INV_X1    g177(.A(G237), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n254), .A3(G214), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(G143), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT17), .B1(new_n366), .B2(new_n244), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n244), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n365), .B(new_n205), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G131), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n371), .B2(KEYINPUT17), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n360), .A2(new_n363), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(G113), .B(G122), .Z(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT85), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n229), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n368), .A2(KEYINPUT18), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n203), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n352), .B2(new_n203), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT18), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n366), .B1(new_n382), .B2(new_n244), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n373), .A2(new_n377), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n377), .B1(new_n373), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n188), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G475), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT19), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n379), .A2(KEYINPUT84), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n350), .A2(new_n351), .B1(new_n379), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(new_n390), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n394), .A2(G146), .B1(new_n368), .B2(new_n370), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n354), .A2(KEYINPUT72), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n358), .A2(new_n397), .A3(G146), .A4(new_n347), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n384), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n376), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT86), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n403), .B(new_n376), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n385), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n389), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n408), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT88), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n210), .A2(G143), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n205), .A2(G128), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n237), .ZN(new_n418));
  XNOR2_X1  g232(.A(G116), .B(G122), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(new_n189), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n189), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT13), .ZN(new_n422));
  OR3_X1    g236(.A1(new_n417), .A2(KEYINPUT89), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n422), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT89), .B1(new_n417), .B2(new_n422), .ZN(new_n425));
  AND4_X1   g239(.A1(new_n416), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  OAI221_X1 g240(.A(new_n418), .B1(new_n420), .B2(new_n421), .C1(new_n426), .C2(new_n237), .ZN(new_n427));
  INV_X1    g241(.A(G116), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n428), .B2(G122), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n419), .B1(KEYINPUT14), .B2(new_n189), .ZN(new_n431));
  INV_X1    g245(.A(new_n418), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n237), .B1(new_n416), .B2(new_n417), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n340), .A2(G217), .A3(new_n254), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT90), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n188), .ZN(new_n439));
  INV_X1    g253(.A(G478), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT15), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n410), .A2(new_n415), .A3(new_n443), .ZN(new_n444));
  NOR4_X1   g258(.A1(new_n288), .A2(new_n338), .A3(new_n342), .A4(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT30), .ZN(new_n447));
  INV_X1    g261(.A(new_n239), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n237), .A2(G137), .ZN(new_n449));
  OAI21_X1  g263(.A(G131), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(new_n245), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n265), .A2(new_n451), .B1(new_n246), .B2(new_n214), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n265), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n246), .A2(new_n214), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n300), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n364), .A2(new_n254), .A3(G210), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT27), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT26), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n463), .B(G101), .Z(new_n464));
  NAND2_X1  g278(.A1(new_n452), .A2(new_n299), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT31), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n457), .A2(new_n300), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n459), .B2(new_n300), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT31), .A3(new_n464), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n452), .A2(new_n299), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT28), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n464), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n468), .A2(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(G472), .A2(G902), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT66), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n446), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n476), .ZN(new_n482));
  INV_X1    g296(.A(new_n471), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT31), .B1(new_n470), .B2(new_n464), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n480), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n473), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n488), .A2(KEYINPUT29), .A3(new_n464), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n464), .A2(new_n473), .A3(new_n475), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n492), .B(new_n493), .C1(new_n470), .C2(new_n464), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n494), .A3(new_n188), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G472), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n481), .A2(new_n487), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G217), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(G234), .B2(new_n188), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT22), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(G137), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n380), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n509));
  OAI211_X1 g323(.A(G119), .B(new_n210), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n506), .A2(new_n507), .B1(new_n304), .B2(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n304), .A2(G128), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G110), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n515), .A2(new_n516), .B1(G119), .B2(new_n210), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT24), .B(G110), .Z(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  AOI211_X1 g334(.A(new_n505), .B(new_n520), .C1(new_n396), .C2(new_n398), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(G110), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n355), .C2(new_n359), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n504), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n520), .B1(new_n396), .B2(new_n398), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n380), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n524), .A3(new_n503), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n529), .A3(new_n188), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n500), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n526), .ZN(new_n535));
  INV_X1    g349(.A(new_n529), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n499), .A2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n497), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n445), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT91), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(new_n216), .Z(G3));
  NAND2_X1  g358(.A1(new_n287), .A2(G469), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n273), .A2(new_n274), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT79), .B1(new_n282), .B2(new_n187), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n342), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n485), .A2(new_n188), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n485), .A2(new_n486), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n553), .A2(new_n534), .A3(new_n539), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n275), .A2(new_n283), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n342), .B1(new_n558), .B2(new_n545), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT92), .A3(new_n554), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n324), .A2(new_n326), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n316), .A2(new_n188), .A3(new_n327), .A4(new_n323), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n562), .A2(new_n337), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n410), .A2(new_n415), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n438), .B(KEYINPUT33), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(G478), .A3(new_n188), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n439), .A2(new_n440), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n564), .A2(new_n336), .A3(new_n565), .A4(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n561), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT34), .B(G104), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G6));
  NAND2_X1  g388(.A1(new_n564), .A2(new_n336), .ZN(new_n575));
  INV_X1    g389(.A(new_n412), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n405), .A2(new_n408), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n413), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n442), .A3(new_n389), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n561), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G107), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G9));
  NAND2_X1  g397(.A1(new_n528), .A2(new_n524), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n504), .A2(KEYINPUT36), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n584), .A2(KEYINPUT36), .A3(new_n504), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n587), .A2(new_n588), .A3(new_n538), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n534), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n445), .A2(new_n552), .A3(new_n551), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT37), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(G110), .Z(G12));
  NOR2_X1   g408(.A1(new_n254), .A2(G900), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(G902), .A3(new_n332), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n333), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n578), .A2(new_n442), .A3(new_n389), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n562), .A2(new_n337), .A3(new_n563), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n601), .A2(new_n602), .A3(new_n590), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n548), .A2(new_n603), .A3(new_n497), .A4(new_n549), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT94), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n559), .A2(new_n606), .A3(new_n497), .A4(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G128), .ZN(G30));
  XOR2_X1   g423(.A(new_n600), .B(KEYINPUT39), .Z(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n559), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT40), .Z(new_n613));
  INV_X1    g427(.A(new_n470), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n464), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n469), .A2(new_n472), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n615), .B1(new_n617), .B2(new_n464), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n619), .B2(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n481), .A3(new_n487), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT98), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n331), .B(KEYINPUT95), .Z(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n565), .A2(new_n442), .ZN(new_n629));
  INV_X1    g443(.A(new_n337), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n590), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n613), .A2(new_n624), .A3(new_n628), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G143), .ZN(G45));
  AND3_X1   g449(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n576), .B1(new_n405), .B2(new_n408), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n636), .A2(new_n637), .A3(new_n406), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n389), .A2(new_n409), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n569), .B(new_n600), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n565), .A2(new_n642), .A3(new_n569), .A4(new_n600), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n564), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n548), .A2(new_n497), .A3(new_n549), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(KEYINPUT101), .A3(new_n564), .A4(new_n643), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n646), .A2(new_n591), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  OR2_X1    g464(.A1(new_n282), .A2(new_n187), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n558), .A2(new_n549), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n652), .A2(new_n571), .A3(new_n653), .A4(new_n541), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n541), .A2(new_n558), .A3(new_n549), .A4(new_n651), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT102), .B1(new_n655), .B2(new_n570), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT41), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G113), .ZN(G15));
  INV_X1    g473(.A(new_n655), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n580), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  NAND4_X1  g476(.A1(new_n558), .A2(new_n549), .A3(new_n564), .A4(new_n651), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n444), .A2(new_n590), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n497), .A3(new_n336), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G119), .ZN(G21));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n540), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT104), .B1(new_n534), .B2(new_n539), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n488), .A2(new_n490), .ZN(new_n671));
  OAI22_X1  g485(.A1(new_n671), .A2(new_n464), .B1(new_n483), .B2(new_n484), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n480), .B(KEYINPUT103), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n550), .A2(G472), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT105), .A4(new_n674), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n575), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n558), .A2(new_n651), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n680), .A2(new_n342), .A3(new_n629), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT106), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n652), .A2(new_n564), .A3(new_n641), .A4(new_n643), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n591), .A2(new_n674), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n641), .A2(new_n643), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n663), .ZN(new_n690));
  INV_X1    g504(.A(new_n687), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(KEYINPUT107), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n285), .B2(new_n256), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n278), .A2(new_n252), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n259), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n284), .A3(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n700), .A2(new_n188), .ZN(new_n701));
  OAI22_X1  g515(.A1(new_n546), .A2(new_n547), .B1(new_n187), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n695), .B1(new_n702), .B2(new_n549), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n187), .B1(new_n700), .B2(new_n188), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n275), .B2(new_n283), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(KEYINPUT109), .A3(new_n342), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n331), .A2(new_n630), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n641), .A2(new_n643), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(KEYINPUT42), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n669), .A2(new_n670), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n497), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT110), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n702), .A2(new_n695), .A3(new_n549), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT109), .B1(new_n705), .B2(new_n342), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n709), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n541), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  INV_X1    g534(.A(new_n712), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n716), .A2(new_n720), .A3(KEYINPUT42), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n713), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  AND2_X1   g538(.A1(new_n541), .A2(new_n708), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n601), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n707), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  NOR2_X1   g543(.A1(new_n638), .A2(new_n639), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n730), .B2(new_n569), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(KEYINPUT43), .A3(new_n569), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT112), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n730), .A2(new_n736), .A3(KEYINPUT43), .A4(new_n569), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n553), .B(new_n591), .C1(new_n733), .C2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n708), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n700), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n286), .A2(new_n744), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(G469), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n558), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n549), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n610), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n739), .A2(KEYINPUT113), .A3(new_n740), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT113), .B1(new_n739), .B2(new_n740), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n743), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  XNOR2_X1  g573(.A(new_n754), .B(KEYINPUT47), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n760), .A2(new_n689), .A3(new_n742), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n497), .A2(new_n540), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n731), .A2(KEYINPUT111), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n731), .A2(KEYINPUT111), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(new_n767), .B1(new_n735), .B2(new_n737), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n765), .B1(new_n768), .B2(new_n333), .ZN(new_n769));
  INV_X1    g583(.A(new_n333), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT118), .B(new_n770), .C1(new_n733), .C2(new_n738), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n677), .A2(new_n678), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n652), .A2(new_n630), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT119), .B1(new_n628), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n625), .B(new_n626), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n630), .A4(new_n652), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n772), .A2(new_n773), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n769), .A2(new_n771), .B1(new_n678), .B2(new_n677), .ZN(new_n782));
  INV_X1    g596(.A(new_n780), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n775), .A4(new_n778), .ZN(new_n784));
  NAND2_X1  g598(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n680), .A2(new_n742), .A3(new_n342), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n772), .A2(new_n691), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n624), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n540), .A3(new_n770), .A4(new_n787), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n565), .A3(new_n569), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n558), .A2(new_n342), .A3(new_n651), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n742), .B1(new_n760), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n793), .B2(new_n782), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n786), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n788), .A4(new_n794), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n772), .A2(new_n721), .A3(new_n787), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT48), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT48), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n800), .A2(new_n801), .B1(new_n664), .B2(new_n782), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n707), .A2(new_n804), .A3(new_n691), .A4(new_n709), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n709), .A2(new_n714), .A3(new_n691), .A4(new_n715), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n591), .A2(new_n389), .A3(new_n578), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n443), .A2(new_n600), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n647), .A2(new_n708), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n807), .A3(new_n728), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  INV_X1    g626(.A(new_n338), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n565), .A2(new_n443), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n557), .A2(new_n813), .A3(new_n560), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n592), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n592), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n654), .A2(new_n656), .B1(new_n445), .B2(new_n541), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n565), .A2(new_n569), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n557), .A2(new_n813), .A3(new_n560), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n679), .A2(new_n681), .B1(new_n660), .B2(new_n580), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n666), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n812), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(KEYINPUT115), .A2(new_n806), .B1(new_n727), .B2(new_n707), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n810), .A4(new_n805), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n723), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT107), .B1(new_n690), .B2(new_n691), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n689), .A2(new_n663), .A3(new_n685), .A4(new_n687), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n608), .B(new_n649), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n705), .A2(new_n342), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n631), .A2(new_n562), .A3(new_n563), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n590), .A2(new_n600), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n624), .A2(new_n838), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT52), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n559), .A2(new_n497), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n645), .B2(new_n644), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n648), .A2(new_n591), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n846), .A2(new_n847), .B1(new_n605), .B2(new_n607), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n693), .A3(new_n849), .A4(new_n842), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n834), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n844), .A2(new_n834), .A3(new_n850), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n832), .B(new_n833), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n825), .B1(new_n818), .B2(new_n819), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n723), .A3(new_n830), .A4(new_n812), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n844), .A2(new_n850), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT53), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n565), .A2(new_n569), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n790), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n833), .B1(new_n855), .B2(new_n856), .ZN(new_n863));
  INV_X1    g677(.A(new_n831), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n812), .A2(new_n820), .A3(new_n826), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n864), .B(new_n865), .C1(new_n852), .C2(new_n851), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n866), .B2(new_n833), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT54), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n803), .A2(new_n860), .A3(new_n862), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n870));
  OAI211_X1 g684(.A(G952), .B(new_n254), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(G953), .B1(new_n869), .B2(KEYINPUT121), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n730), .A2(new_n549), .A3(new_n569), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n711), .A2(new_n337), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n873), .B(new_n874), .C1(KEYINPUT49), .C2(new_n680), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n680), .A2(KEYINPUT49), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n776), .A3(new_n789), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n872), .A3(new_n877), .ZN(G75));
  NAND4_X1  g692(.A1(new_n853), .A2(G210), .A3(G902), .A4(new_n857), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n294), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT55), .Z(new_n884));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  INV_X1    g700(.A(new_n884), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n886), .B(new_n887), .C1(new_n879), .C2(new_n880), .ZN(new_n888));
  OAI211_X1 g702(.A(G902), .B(new_n857), .C1(new_n866), .C2(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT123), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n853), .A2(new_n891), .A3(G902), .A4(new_n857), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n326), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n880), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n885), .A2(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n254), .A2(G952), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT124), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(G51));
  AND2_X1   g712(.A1(new_n890), .A2(new_n892), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(new_n747), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n858), .B(KEYINPUT54), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n748), .B(KEYINPUT57), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n901), .A2(new_n902), .B1(new_n272), .B2(new_n269), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n896), .B1(new_n900), .B2(new_n903), .ZN(G54));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n890), .B2(new_n892), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n906), .A2(G475), .A3(new_n405), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n405), .B1(new_n906), .B2(G475), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n896), .ZN(G60));
  INV_X1    g723(.A(new_n566), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n860), .A2(new_n868), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n897), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n858), .B(new_n859), .ZN(new_n916));
  INV_X1    g730(.A(new_n913), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n566), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(G63));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  OAI211_X1 g736(.A(new_n857), .B(new_n922), .C1(new_n866), .C2(KEYINPUT53), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n853), .A2(new_n925), .A3(new_n857), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n535), .A2(new_n536), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n915), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n587), .A2(new_n588), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n924), .B2(new_n926), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n920), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n932), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n924), .B(new_n926), .C1(new_n536), .C2(new_n535), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n934), .A2(KEYINPUT61), .A3(new_n935), .A4(new_n915), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(G66));
  AOI21_X1  g751(.A(new_n254), .B1(new_n334), .B2(new_n292), .ZN(new_n938));
  INV_X1    g752(.A(new_n854), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n254), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n882), .B1(G898), .B2(new_n254), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(G69));
  XOR2_X1   g756(.A(new_n459), .B(new_n394), .Z(new_n943));
  INV_X1    g757(.A(new_n837), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n634), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT62), .Z(new_n946));
  INV_X1    g760(.A(new_n612), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n725), .C1(new_n822), .C2(new_n814), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n758), .A3(new_n763), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(new_n254), .ZN(new_n950));
  INV_X1    g764(.A(new_n943), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n763), .A2(new_n728), .A3(new_n758), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n755), .A2(new_n721), .A3(new_n839), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n723), .A2(new_n944), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n254), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n595), .B(KEYINPUT127), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(G227), .A2(G900), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n957), .A2(KEYINPUT126), .B1(new_n254), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n958), .B(new_n960), .Z(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n949), .B2(new_n939), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n464), .A3(new_n614), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n614), .A2(new_n464), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n952), .A2(new_n939), .A3(new_n954), .ZN(new_n967));
  INV_X1    g781(.A(new_n963), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n965), .B(new_n969), .C1(G952), .C2(new_n254), .ZN(new_n970));
  INV_X1    g784(.A(new_n966), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n867), .A2(new_n615), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n963), .B2(new_n972), .ZN(G57));
endmodule


