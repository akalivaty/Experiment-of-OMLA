

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732;

  XNOR2_X1 U363 ( .A(n404), .B(n403), .ZN(n670) );
  INV_X1 U364 ( .A(G953), .ZN(n489) );
  AND2_X2 U365 ( .A1(n363), .A2(n360), .ZN(n359) );
  AND2_X2 U366 ( .A1(n398), .A2(n397), .ZN(n396) );
  AND2_X4 U367 ( .A1(n602), .A2(n601), .ZN(n700) );
  XNOR2_X2 U368 ( .A(n715), .B(n430), .ZN(n621) );
  XNOR2_X2 U369 ( .A(n491), .B(n414), .ZN(n691) );
  XNOR2_X2 U370 ( .A(n721), .B(n481), .ZN(n491) );
  NOR2_X2 U371 ( .A1(n691), .A2(G902), .ZN(n494) );
  XNOR2_X1 U372 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n423) );
  XOR2_X1 U373 ( .A(KEYINPUT90), .B(KEYINPUT78), .Z(n424) );
  OR2_X1 U374 ( .A1(n540), .A2(n662), .ZN(n355) );
  XNOR2_X1 U375 ( .A(n514), .B(n488), .ZN(n573) );
  XOR2_X1 U376 ( .A(KEYINPUT59), .B(n695), .Z(n696) );
  XNOR2_X1 U377 ( .A(n424), .B(n423), .ZN(n427) );
  XNOR2_X1 U378 ( .A(n401), .B(G143), .ZN(n462) );
  XNOR2_X2 U379 ( .A(n577), .B(n437), .ZN(n581) );
  XNOR2_X2 U380 ( .A(n511), .B(n510), .ZN(n730) );
  XNOR2_X2 U381 ( .A(n421), .B(n485), .ZN(n715) );
  XNOR2_X1 U382 ( .A(n536), .B(n372), .ZN(n353) );
  NAND2_X1 U383 ( .A1(n541), .A2(n355), .ZN(n354) );
  INV_X1 U384 ( .A(KEYINPUT106), .ZN(n372) );
  XNOR2_X1 U385 ( .A(n479), .B(n384), .ZN(n721) );
  XNOR2_X1 U386 ( .A(n480), .B(n385), .ZN(n384) );
  XNOR2_X1 U387 ( .A(n386), .B(KEYINPUT4), .ZN(n385) );
  INV_X1 U388 ( .A(G137), .ZN(n386) );
  OR2_X1 U389 ( .A1(n609), .A2(G902), .ZN(n404) );
  XNOR2_X1 U390 ( .A(n418), .B(G101), .ZN(n382) );
  INV_X1 U391 ( .A(G146), .ZN(n481) );
  NAND2_X1 U392 ( .A1(n521), .A2(n682), .ZN(n377) );
  INV_X1 U393 ( .A(KEYINPUT22), .ZN(n373) );
  XNOR2_X1 U394 ( .A(n367), .B(n590), .ZN(n402) );
  NAND2_X1 U395 ( .A1(n340), .A2(n348), .ZN(n367) );
  XNOR2_X1 U396 ( .A(KEYINPUT15), .B(G902), .ZN(n598) );
  OR2_X1 U397 ( .A1(n654), .A2(KEYINPUT87), .ZN(n397) );
  XNOR2_X1 U398 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n496) );
  XNOR2_X1 U399 ( .A(G128), .B(KEYINPUT75), .ZN(n498) );
  XNOR2_X1 U400 ( .A(n462), .B(n461), .ZN(n479) );
  INV_X1 U401 ( .A(G134), .ZN(n461) );
  XNOR2_X1 U402 ( .A(G122), .B(G116), .ZN(n463) );
  XOR2_X1 U403 ( .A(KEYINPUT102), .B(G107), .Z(n464) );
  XNOR2_X1 U404 ( .A(n379), .B(n378), .ZN(n495) );
  INV_X1 U405 ( .A(KEYINPUT8), .ZN(n378) );
  NAND2_X1 U406 ( .A1(n489), .A2(G234), .ZN(n379) );
  INV_X1 U407 ( .A(KEYINPUT10), .ZN(n450) );
  INV_X1 U408 ( .A(n573), .ZN(n407) );
  XNOR2_X1 U409 ( .A(n558), .B(KEYINPUT39), .ZN(n597) );
  INV_X1 U410 ( .A(KEYINPUT34), .ZN(n390) );
  INV_X1 U411 ( .A(n513), .ZN(n403) );
  INV_X1 U412 ( .A(KEYINPUT0), .ZN(n444) );
  OR2_X1 U413 ( .A1(n701), .A2(G902), .ZN(n509) );
  XNOR2_X1 U414 ( .A(n492), .B(G101), .ZN(n414) );
  XNOR2_X1 U415 ( .A(n490), .B(n392), .ZN(n391) );
  INV_X1 U416 ( .A(KEYINPUT70), .ZN(n365) );
  INV_X1 U417 ( .A(KEYINPUT44), .ZN(n361) );
  XNOR2_X1 U418 ( .A(G119), .B(G110), .ZN(n500) );
  XNOR2_X1 U419 ( .A(KEYINPUT24), .B(G137), .ZN(n499) );
  XNOR2_X1 U420 ( .A(KEYINPUT77), .B(KEYINPUT89), .ZN(n425) );
  XNOR2_X1 U421 ( .A(n422), .B(n400), .ZN(n399) );
  INV_X1 U422 ( .A(KEYINPUT4), .ZN(n400) );
  NAND2_X1 U423 ( .A1(n375), .A2(n661), .ZN(n672) );
  XNOR2_X1 U424 ( .A(n513), .B(n487), .ZN(n488) );
  AND2_X1 U425 ( .A1(n402), .A2(n345), .ZN(n722) );
  XNOR2_X1 U426 ( .A(n387), .B(G131), .ZN(n480) );
  INV_X1 U427 ( .A(KEYINPUT66), .ZN(n387) );
  XNOR2_X1 U428 ( .A(G143), .B(G122), .ZN(n453) );
  XOR2_X1 U429 ( .A(G104), .B(G113), .Z(n454) );
  NAND2_X1 U430 ( .A1(n350), .A2(n413), .ZN(n412) );
  NAND2_X1 U431 ( .A1(n598), .A2(KEYINPUT83), .ZN(n413) );
  XNOR2_X1 U432 ( .A(G140), .B(KEYINPUT76), .ZN(n392) );
  NAND2_X1 U433 ( .A1(n395), .A2(n394), .ZN(n393) );
  AND2_X1 U434 ( .A1(n654), .A2(KEYINPUT87), .ZN(n394) );
  XNOR2_X1 U435 ( .A(n491), .B(n405), .ZN(n609) );
  XNOR2_X1 U436 ( .A(n486), .B(n343), .ZN(n405) );
  XNOR2_X1 U437 ( .A(n357), .B(n417), .ZN(n421) );
  XNOR2_X1 U438 ( .A(n416), .B(G122), .ZN(n417) );
  INV_X1 U439 ( .A(KEYINPUT16), .ZN(n416) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n701) );
  XNOR2_X1 U441 ( .A(n503), .B(n497), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n719), .B(n496), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n479), .B(n471), .ZN(n603) );
  XNOR2_X1 U444 ( .A(n560), .B(n559), .ZN(n617) );
  INV_X1 U445 ( .A(n584), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n377), .B(n390), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n528), .B(n527), .ZN(n642) );
  INV_X1 U448 ( .A(KEYINPUT31), .ZN(n527) );
  INV_X1 U449 ( .A(n592), .ZN(n512) );
  INV_X1 U450 ( .A(n550), .ZN(n371) );
  XNOR2_X1 U451 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U452 ( .A(KEYINPUT46), .B(n571), .ZN(n340) );
  NOR2_X1 U453 ( .A1(KEYINPUT83), .A2(n598), .ZN(n341) );
  INV_X1 U454 ( .A(n663), .ZN(n368) );
  XOR2_X1 U455 ( .A(n370), .B(KEYINPUT107), .Z(n342) );
  XOR2_X1 U456 ( .A(n482), .B(KEYINPUT5), .Z(n343) );
  OR2_X1 U457 ( .A1(G902), .A2(n603), .ZN(n344) );
  AND2_X1 U458 ( .A1(n647), .A2(n614), .ZN(n345) );
  AND2_X1 U459 ( .A1(n706), .A2(n409), .ZN(n346) );
  OR2_X1 U460 ( .A1(n519), .A2(n518), .ZN(n347) );
  AND2_X1 U461 ( .A1(n589), .A2(n588), .ZN(n348) );
  AND2_X1 U462 ( .A1(n345), .A2(n341), .ZN(n349) );
  NAND2_X1 U463 ( .A1(n599), .A2(KEYINPUT2), .ZN(n350) );
  XOR2_X1 U464 ( .A(n609), .B(KEYINPUT62), .Z(n351) );
  NAND2_X1 U465 ( .A1(n359), .A2(n358), .ZN(n520) );
  AND2_X1 U466 ( .A1(n362), .A2(n361), .ZN(n360) );
  INV_X1 U467 ( .A(n355), .ZN(n616) );
  XNOR2_X1 U468 ( .A(n352), .B(KEYINPUT86), .ZN(n542) );
  NOR2_X2 U469 ( .A1(n354), .A2(n353), .ZN(n352) );
  NAND2_X1 U470 ( .A1(n356), .A2(n512), .ZN(n516) );
  NAND2_X1 U471 ( .A1(n356), .A2(n573), .ZN(n538) );
  XNOR2_X2 U472 ( .A(n374), .B(n373), .ZN(n356) );
  XNOR2_X1 U473 ( .A(n357), .B(n391), .ZN(n492) );
  XNOR2_X2 U474 ( .A(n415), .B(G110), .ZN(n357) );
  NAND2_X1 U475 ( .A1(n519), .A2(n365), .ZN(n358) );
  NAND2_X1 U476 ( .A1(n618), .A2(n365), .ZN(n362) );
  NAND2_X1 U477 ( .A1(n366), .A2(n364), .ZN(n363) );
  NOR2_X1 U478 ( .A1(n618), .A2(n365), .ZN(n364) );
  INV_X1 U479 ( .A(n519), .ZN(n366) );
  NAND2_X1 U480 ( .A1(n730), .A2(n615), .ZN(n519) );
  NOR2_X1 U481 ( .A1(n346), .A2(n412), .ZN(n411) );
  NAND2_X1 U482 ( .A1(n369), .A2(n368), .ZN(n517) );
  INV_X1 U483 ( .A(n662), .ZN(n369) );
  NOR2_X1 U484 ( .A1(n617), .A2(n732), .ZN(n571) );
  NAND2_X1 U485 ( .A1(n411), .A2(n410), .ZN(n602) );
  XNOR2_X1 U486 ( .A(n462), .B(n399), .ZN(n429) );
  XNOR2_X2 U487 ( .A(n544), .B(KEYINPUT45), .ZN(n706) );
  NAND2_X1 U488 ( .A1(n618), .A2(KEYINPUT44), .ZN(n541) );
  INV_X1 U489 ( .A(n404), .ZN(n514) );
  XNOR2_X2 U490 ( .A(n522), .B(KEYINPUT1), .ZN(n537) );
  NAND2_X1 U491 ( .A1(n579), .A2(n662), .ZN(n370) );
  INV_X1 U492 ( .A(n521), .ZN(n525) );
  AND2_X1 U493 ( .A1(n521), .A2(n371), .ZN(n523) );
  XNOR2_X2 U494 ( .A(n445), .B(n444), .ZN(n521) );
  NAND2_X1 U495 ( .A1(n521), .A2(n478), .ZN(n374) );
  NOR2_X1 U496 ( .A1(n525), .A2(n375), .ZN(n526) );
  INV_X1 U497 ( .A(n408), .ZN(n375) );
  AND2_X2 U498 ( .A1(n665), .A2(n537), .ZN(n408) );
  NAND2_X1 U499 ( .A1(n376), .A2(n389), .ZN(n388) );
  XNOR2_X2 U500 ( .A(n406), .B(KEYINPUT33), .ZN(n682) );
  XNOR2_X2 U501 ( .A(n383), .B(n382), .ZN(n485) );
  XNOR2_X2 U502 ( .A(n420), .B(n419), .ZN(n383) );
  XNOR2_X2 U503 ( .A(n388), .B(KEYINPUT35), .ZN(n618) );
  NAND2_X2 U504 ( .A1(n396), .A2(n393), .ZN(n577) );
  INV_X1 U505 ( .A(n555), .ZN(n395) );
  NAND2_X1 U506 ( .A1(n555), .A2(n436), .ZN(n398) );
  XNOR2_X2 U507 ( .A(G128), .B(KEYINPUT79), .ZN(n401) );
  XNOR2_X2 U508 ( .A(n509), .B(n508), .ZN(n662) );
  AND2_X1 U509 ( .A1(n402), .A2(n349), .ZN(n409) );
  NAND2_X1 U510 ( .A1(n408), .A2(n407), .ZN(n406) );
  NAND2_X1 U511 ( .A1(n706), .A2(n722), .ZN(n648) );
  NAND2_X1 U512 ( .A1(n648), .A2(KEYINPUT83), .ZN(n410) );
  XNOR2_X1 U513 ( .A(n610), .B(n351), .ZN(n612) );
  BUF_X1 U514 ( .A(n522), .Z(n564) );
  AND2_X1 U515 ( .A1(n567), .A2(n368), .ZN(n478) );
  BUF_X1 U516 ( .A(n537), .Z(n592) );
  INV_X1 U517 ( .A(n703), .ZN(n611) );
  XNOR2_X2 U518 ( .A(G107), .B(G104), .ZN(n415) );
  XNOR2_X2 U519 ( .A(G113), .B(KEYINPUT3), .ZN(n419) );
  INV_X1 U520 ( .A(KEYINPUT68), .ZN(n418) );
  XNOR2_X2 U521 ( .A(G116), .B(G119), .ZN(n420) );
  NAND2_X1 U522 ( .A1(G224), .A2(n489), .ZN(n422) );
  XNOR2_X2 U523 ( .A(G146), .B(G125), .ZN(n452) );
  XNOR2_X1 U524 ( .A(n425), .B(n452), .ZN(n426) );
  XNOR2_X1 U525 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U526 ( .A(n428), .B(n429), .ZN(n430) );
  NAND2_X1 U527 ( .A1(n621), .A2(n598), .ZN(n434) );
  XOR2_X1 U528 ( .A(KEYINPUT91), .B(KEYINPUT80), .Z(n432) );
  OR2_X1 U529 ( .A1(G902), .A2(G237), .ZN(n435) );
  NAND2_X1 U530 ( .A1(G210), .A2(n435), .ZN(n431) );
  XNOR2_X1 U531 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X2 U532 ( .A(n434), .B(n433), .ZN(n555) );
  NAND2_X1 U533 ( .A1(G214), .A2(n435), .ZN(n654) );
  INV_X1 U534 ( .A(KEYINPUT87), .ZN(n436) );
  XNOR2_X1 U535 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n437) );
  NAND2_X1 U536 ( .A1(G237), .A2(G234), .ZN(n438) );
  XNOR2_X1 U537 ( .A(n438), .B(KEYINPUT14), .ZN(n439) );
  XNOR2_X1 U538 ( .A(KEYINPUT72), .B(n439), .ZN(n440) );
  NAND2_X1 U539 ( .A1(G952), .A2(n440), .ZN(n680) );
  NOR2_X1 U540 ( .A1(G953), .A2(n680), .ZN(n548) );
  AND2_X1 U541 ( .A1(n440), .A2(G902), .ZN(n545) );
  NOR2_X1 U542 ( .A1(G898), .A2(n489), .ZN(n716) );
  NAND2_X1 U543 ( .A1(n545), .A2(n716), .ZN(n441) );
  XOR2_X1 U544 ( .A(KEYINPUT92), .B(n441), .Z(n442) );
  OR2_X1 U545 ( .A1(n548), .A2(n442), .ZN(n443) );
  NAND2_X1 U546 ( .A1(n581), .A2(n443), .ZN(n445) );
  XNOR2_X1 U547 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n459) );
  XNOR2_X1 U548 ( .A(n480), .B(KEYINPUT12), .ZN(n449) );
  XOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n447) );
  NOR2_X1 U550 ( .A1(G953), .A2(G237), .ZN(n483) );
  NAND2_X1 U551 ( .A1(n483), .A2(G214), .ZN(n446) );
  XNOR2_X1 U552 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U553 ( .A(n449), .B(n448), .ZN(n457) );
  XNOR2_X1 U554 ( .A(n450), .B(G140), .ZN(n451) );
  XNOR2_X1 U555 ( .A(n451), .B(n452), .ZN(n719) );
  XNOR2_X1 U556 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n719), .B(n455), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n695) );
  NOR2_X1 U559 ( .A1(G902), .A2(n695), .ZN(n458) );
  XNOR2_X1 U560 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U561 ( .A(n460), .B(G475), .ZN(n529) );
  XNOR2_X1 U562 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U563 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n466) );
  XNOR2_X1 U564 ( .A(KEYINPUT103), .B(KEYINPUT9), .ZN(n465) );
  XNOR2_X1 U565 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U566 ( .A(n468), .B(n467), .Z(n470) );
  NAND2_X1 U567 ( .A1(G217), .A2(n495), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U569 ( .A(G478), .B(n344), .ZN(n532) );
  NOR2_X1 U570 ( .A1(n529), .A2(n532), .ZN(n567) );
  NAND2_X1 U571 ( .A1(n598), .A2(G234), .ZN(n473) );
  INV_X1 U572 ( .A(KEYINPUT20), .ZN(n472) );
  XNOR2_X1 U573 ( .A(n473), .B(n472), .ZN(n504) );
  INV_X1 U574 ( .A(G221), .ZN(n474) );
  OR2_X1 U575 ( .A1(n504), .A2(n474), .ZN(n477) );
  INV_X1 U576 ( .A(KEYINPUT95), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n475), .B(KEYINPUT21), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n477), .B(n476), .ZN(n663) );
  XNOR2_X1 U579 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n482) );
  NAND2_X1 U580 ( .A1(n483), .A2(G210), .ZN(n484) );
  XNOR2_X1 U581 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U582 ( .A(KEYINPUT71), .B(G472), .Z(n513) );
  INV_X1 U583 ( .A(KEYINPUT6), .ZN(n487) );
  NAND2_X1 U584 ( .A1(G227), .A2(n489), .ZN(n490) );
  INV_X1 U585 ( .A(G469), .ZN(n493) );
  XNOR2_X2 U586 ( .A(n494), .B(n493), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n537), .B(KEYINPUT88), .ZN(n579) );
  NAND2_X1 U588 ( .A1(n495), .A2(G221), .ZN(n497) );
  XNOR2_X1 U589 ( .A(n499), .B(n498), .ZN(n502) );
  XNOR2_X1 U590 ( .A(n500), .B(KEYINPUT69), .ZN(n501) );
  XNOR2_X1 U591 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U592 ( .A(n504), .ZN(n505) );
  NAND2_X1 U593 ( .A1(n505), .A2(G217), .ZN(n507) );
  XNOR2_X1 U594 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n506) );
  XNOR2_X1 U595 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X2 U596 ( .A1(n538), .A2(n342), .ZN(n511) );
  XOR2_X1 U597 ( .A(KEYINPUT64), .B(KEYINPUT32), .Z(n510) );
  NAND2_X1 U598 ( .A1(n670), .A2(n662), .ZN(n515) );
  OR2_X1 U599 ( .A1(n516), .A2(n515), .ZN(n615) );
  XNOR2_X1 U600 ( .A(n517), .B(KEYINPUT65), .ZN(n665) );
  NAND2_X1 U601 ( .A1(n529), .A2(n532), .ZN(n584) );
  NAND2_X1 U602 ( .A1(KEYINPUT70), .A2(KEYINPUT44), .ZN(n518) );
  NAND2_X1 U603 ( .A1(n520), .A2(n347), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n564), .A2(n665), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n523), .B(KEYINPUT96), .ZN(n524) );
  NAND2_X1 U606 ( .A1(n524), .A2(n670), .ZN(n629) );
  INV_X1 U607 ( .A(n670), .ZN(n661) );
  NAND2_X1 U608 ( .A1(n526), .A2(n661), .ZN(n528) );
  NAND2_X1 U609 ( .A1(n629), .A2(n642), .ZN(n535) );
  XNOR2_X1 U610 ( .A(n529), .B(KEYINPUT101), .ZN(n533) );
  OR2_X1 U611 ( .A1(n533), .A2(n532), .ZN(n531) );
  INV_X1 U612 ( .A(KEYINPUT105), .ZN(n530) );
  XNOR2_X1 U613 ( .A(n531), .B(n530), .ZN(n640) );
  NAND2_X1 U614 ( .A1(n533), .A2(n532), .ZN(n643) );
  AND2_X1 U615 ( .A1(n640), .A2(n643), .ZN(n651) );
  INV_X1 U616 ( .A(n651), .ZN(n534) );
  NAND2_X1 U617 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U618 ( .A1(n538), .A2(n592), .ZN(n539) );
  XNOR2_X1 U619 ( .A(n539), .B(KEYINPUT85), .ZN(n540) );
  NAND2_X1 U620 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U621 ( .A1(G953), .A2(n545), .ZN(n546) );
  NOR2_X1 U622 ( .A1(G900), .A2(n546), .ZN(n547) );
  OR2_X1 U623 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U624 ( .A(n549), .B(KEYINPUT81), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n550), .A2(n561), .ZN(n554) );
  INV_X1 U626 ( .A(n654), .ZN(n551) );
  NOR2_X1 U627 ( .A1(n670), .A2(n551), .ZN(n552) );
  XNOR2_X1 U628 ( .A(n552), .B(KEYINPUT30), .ZN(n553) );
  AND2_X1 U629 ( .A1(n554), .A2(n553), .ZN(n586) );
  BUF_X1 U630 ( .A(n555), .Z(n556) );
  XOR2_X1 U631 ( .A(KEYINPUT73), .B(KEYINPUT38), .Z(n557) );
  XNOR2_X1 U632 ( .A(n556), .B(n557), .ZN(n653) );
  NAND2_X1 U633 ( .A1(n586), .A2(n653), .ZN(n558) );
  INV_X1 U634 ( .A(n640), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n597), .A2(n575), .ZN(n560) );
  XOR2_X1 U636 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n559) );
  NOR2_X1 U637 ( .A1(n561), .A2(n663), .ZN(n562) );
  NAND2_X1 U638 ( .A1(n562), .A2(n662), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n670), .A2(n572), .ZN(n563) );
  XOR2_X1 U640 ( .A(KEYINPUT28), .B(n563), .Z(n566) );
  XNOR2_X1 U641 ( .A(n564), .B(KEYINPUT109), .ZN(n565) );
  NOR2_X1 U642 ( .A1(n566), .A2(n565), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n654), .A2(n653), .ZN(n650) );
  INV_X1 U644 ( .A(n567), .ZN(n656) );
  NOR2_X1 U645 ( .A1(n650), .A2(n656), .ZN(n569) );
  XNOR2_X1 U646 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n568) );
  XNOR2_X1 U647 ( .A(n569), .B(n568), .ZN(n681) );
  NAND2_X1 U648 ( .A1(n582), .A2(n681), .ZN(n570) );
  XOR2_X1 U649 ( .A(n570), .B(KEYINPUT42), .Z(n732) );
  NOR2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(n574), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n591) );
  NOR2_X1 U653 ( .A1(n577), .A2(n591), .ZN(n578) );
  XNOR2_X1 U654 ( .A(KEYINPUT36), .B(n578), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n646) );
  XNOR2_X1 U656 ( .A(n646), .B(KEYINPUT84), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n638) );
  NOR2_X1 U658 ( .A1(n638), .A2(n651), .ZN(n583) );
  XOR2_X1 U659 ( .A(n583), .B(KEYINPUT47), .Z(n587) );
  NOR2_X1 U660 ( .A1(n556), .A2(n584), .ZN(n585) );
  AND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n637) );
  NOR2_X1 U662 ( .A1(n587), .A2(n637), .ZN(n588) );
  XNOR2_X1 U663 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n593), .A2(n654), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT43), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n595), .A2(n556), .ZN(n647) );
  INV_X1 U668 ( .A(n643), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n614) );
  INV_X1 U670 ( .A(n598), .ZN(n599) );
  INV_X1 U671 ( .A(n648), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n600), .A2(KEYINPUT2), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n700), .A2(G478), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(n606) );
  INV_X1 U675 ( .A(G952), .ZN(n605) );
  AND2_X1 U676 ( .A1(n605), .A2(G953), .ZN(n703) );
  NOR2_X2 U677 ( .A1(n606), .A2(n703), .ZN(n608) );
  INV_X1 U678 ( .A(KEYINPUT119), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(G63) );
  NAND2_X1 U680 ( .A1(n700), .A2(G472), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U683 ( .A(n614), .B(G134), .ZN(G36) );
  XNOR2_X1 U684 ( .A(n615), .B(G110), .ZN(G12) );
  XOR2_X1 U685 ( .A(G101), .B(n616), .Z(G3) );
  XOR2_X1 U686 ( .A(G131), .B(n617), .Z(G33) );
  XNOR2_X1 U687 ( .A(G122), .B(KEYINPUT126), .ZN(n619) );
  XOR2_X1 U688 ( .A(n619), .B(n618), .Z(G24) );
  NAND2_X1 U689 ( .A1(n700), .A2(G210), .ZN(n623) );
  XOR2_X1 U690 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n624), .A2(n611), .ZN(n626) );
  INV_X1 U694 ( .A(KEYINPUT56), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(G51) );
  NOR2_X1 U696 ( .A1(n640), .A2(n629), .ZN(n627) );
  XOR2_X1 U697 ( .A(KEYINPUT112), .B(n627), .Z(n628) );
  XNOR2_X1 U698 ( .A(G104), .B(n628), .ZN(G6) );
  NOR2_X1 U699 ( .A1(n643), .A2(n629), .ZN(n634) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n631) );
  XNOR2_X1 U701 ( .A(G107), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(KEYINPUT113), .B(n632), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(G9) );
  NOR2_X1 U705 ( .A1(n643), .A2(n638), .ZN(n636) );
  XNOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(G30) );
  XOR2_X1 U708 ( .A(G143), .B(n637), .Z(G45) );
  NOR2_X1 U709 ( .A1(n640), .A2(n638), .ZN(n639) );
  XOR2_X1 U710 ( .A(G146), .B(n639), .Z(G48) );
  NOR2_X1 U711 ( .A1(n640), .A2(n642), .ZN(n641) );
  XOR2_X1 U712 ( .A(G113), .B(n641), .Z(G15) );
  NOR2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U714 ( .A(G116), .B(n644), .Z(G18) );
  XOR2_X1 U715 ( .A(G125), .B(KEYINPUT37), .Z(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G27) );
  XNOR2_X1 U717 ( .A(G140), .B(n647), .ZN(G42) );
  NAND2_X1 U718 ( .A1(n648), .A2(KEYINPUT82), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n649), .B(KEYINPUT2), .ZN(n686) );
  NOR2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT116), .B(n652), .Z(n659) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U724 ( .A(KEYINPUT115), .B(n657), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U726 ( .A1(n682), .A2(n660), .ZN(n676) );
  NAND2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U728 ( .A(KEYINPUT49), .B(n664), .Z(n668) );
  NOR2_X1 U729 ( .A1(n665), .A2(n537), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT50), .B(n666), .Z(n667) );
  NAND2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U734 ( .A(KEYINPUT51), .B(n673), .ZN(n674) );
  NAND2_X1 U735 ( .A1(n674), .A2(n681), .ZN(n675) );
  NAND2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U737 ( .A(n677), .B(KEYINPUT117), .ZN(n678) );
  XNOR2_X1 U738 ( .A(n678), .B(KEYINPUT52), .ZN(n679) );
  NOR2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n684) );
  AND2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U743 ( .A1(G953), .A2(n687), .ZN(n689) );
  XNOR2_X1 U744 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n688) );
  XNOR2_X1 U745 ( .A(n689), .B(n688), .ZN(G75) );
  NAND2_X1 U746 ( .A1(n700), .A2(G469), .ZN(n693) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n690) );
  XNOR2_X1 U748 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U749 ( .A1(n703), .A2(n694), .ZN(G54) );
  NAND2_X1 U750 ( .A1(n700), .A2(G475), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X2 U752 ( .A1(n698), .A2(n703), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n699), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U754 ( .A1(n700), .A2(G217), .ZN(n702) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X2 U756 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U757 ( .A(n705), .B(KEYINPUT120), .ZN(G66) );
  INV_X1 U758 ( .A(n706), .ZN(n707) );
  NOR2_X1 U759 ( .A1(n707), .A2(G953), .ZN(n714) );
  XOR2_X1 U760 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n709) );
  NAND2_X1 U761 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U762 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U763 ( .A(KEYINPUT121), .B(n710), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n711), .A2(G898), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n712), .B(KEYINPUT123), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n715), .A2(n716), .ZN(n717) );
  XOR2_X1 U768 ( .A(n718), .B(n717), .Z(G69) );
  XNOR2_X1 U769 ( .A(n719), .B(KEYINPUT124), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n725) );
  XNOR2_X1 U771 ( .A(n722), .B(n725), .ZN(n723) );
  NOR2_X1 U772 ( .A1(n723), .A2(G953), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(KEYINPUT125), .ZN(n729) );
  XNOR2_X1 U774 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U775 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U778 ( .A(G119), .B(KEYINPUT127), .Z(n731) );
  XNOR2_X1 U779 ( .A(n730), .B(n731), .ZN(G21) );
  XOR2_X1 U780 ( .A(G137), .B(n732), .Z(G39) );
endmodule

