//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT91), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n210), .A2(KEYINPUT92), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(KEYINPUT92), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(KEYINPUT16), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n208), .A2(KEYINPUT91), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n208), .A2(KEYINPUT91), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(G1gat), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT93), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n213), .A2(new_n216), .B1(new_n217), .B2(G8gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(G8gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n213), .A2(KEYINPUT93), .A3(new_n222), .A4(new_n216), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G43gat), .B(G50gat), .Z(new_n227));
  INV_X1    g026(.A(KEYINPUT15), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OR3_X1    g030(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT88), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n233), .B2(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(G29gat), .A2(G36gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT89), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n229), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n227), .A2(new_n228), .B1(new_n232), .B2(new_n230), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n229), .A2(new_n239), .A3(new_n237), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n221), .A2(KEYINPUT94), .A3(new_n223), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT95), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n226), .A2(KEYINPUT95), .A3(new_n242), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n241), .A2(KEYINPUT17), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT90), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n241), .A2(KEYINPUT17), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n224), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n248), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n207), .B1(new_n256), .B2(KEYINPUT97), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n248), .A2(KEYINPUT18), .A3(new_n249), .A4(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n226), .A2(new_n243), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n241), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n248), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n249), .B(KEYINPUT13), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n254), .A2(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT97), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n254), .B2(new_n255), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n266), .B(new_n258), .C1(new_n268), .C2(new_n207), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(G169gat), .ZN(new_n274));
  INV_X1    g073(.A(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n280), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT28), .B1(new_n286), .B2(G190gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT69), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n284), .A2(new_n287), .A3(new_n288), .A4(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT23), .ZN(new_n294));
  OAI22_X1  g093(.A1(KEYINPUT66), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n278), .B(new_n294), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(KEYINPUT24), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n299), .A2(new_n307), .A3(KEYINPUT68), .A4(KEYINPUT25), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G190gat), .ZN(new_n310));
  OAI211_X1 g109(.A(KEYINPUT25), .B(new_n301), .C1(new_n310), .C2(new_n300), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n311), .B2(new_n298), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n276), .A3(new_n296), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n317), .A2(KEYINPUT67), .A3(new_n278), .A4(new_n294), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n318), .A3(new_n307), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n293), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n272), .B(new_n273), .C1(new_n322), .C2(KEYINPUT29), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT74), .B1(new_n322), .B2(new_n273), .ZN(new_n324));
  INV_X1    g123(.A(new_n273), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n301), .B1(new_n310), .B2(new_n300), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n314), .B2(new_n298), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT25), .B1(new_n327), .B2(new_n318), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n312), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n292), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n323), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335));
  INV_X1    g134(.A(G211gat), .ZN(new_n336));
  INV_X1    g135(.A(G218gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n334), .A3(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n333), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n273), .C1(new_n322), .C2(KEYINPUT29), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT73), .B1(new_n330), .B2(new_n325), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n332), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n344), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT37), .ZN(new_n354));
  XOR2_X1   g153(.A(G8gat), .B(G36gat), .Z(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT75), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(KEYINPUT37), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n345), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT38), .ZN(new_n362));
  INV_X1    g161(.A(new_n358), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n352), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT2), .ZN(new_n367));
  OR2_X1    g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(G155gat), .B2(G162gat), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n370), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n365), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n370), .A2(new_n373), .ZN(new_n377));
  INV_X1    g176(.A(new_n371), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT3), .A3(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G127gat), .B(G134gat), .Z(new_n382));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(KEYINPUT1), .B2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G113gat), .B(G120gat), .Z(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  XNOR2_X1  g185(.A(G127gat), .B(G134gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n384), .A2(new_n388), .A3(KEYINPUT77), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT77), .B1(new_n384), .B2(new_n388), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n376), .B(new_n381), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n374), .A2(new_n375), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n384), .A2(new_n388), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n395), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n380), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT4), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n391), .A2(new_n392), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n389), .B2(new_n390), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n398), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n392), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n396), .A2(new_n399), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n406), .A2(KEYINPUT5), .A3(new_n392), .A4(new_n391), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT6), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n412), .B(KEYINPUT83), .Z(new_n415));
  NAND3_X1  g214(.A1(new_n405), .A2(new_n415), .A3(new_n407), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT6), .A4(new_n412), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n364), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n351), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n347), .B(new_n420), .C1(new_n332), .C2(new_n348), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n333), .B2(new_n344), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT37), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT38), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n360), .A3(new_n424), .A4(new_n358), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT86), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n419), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n362), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n342), .B2(new_n343), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n394), .B1(new_n430), .B2(KEYINPUT3), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n394), .B(KEYINPUT80), .C1(new_n430), .C2(KEYINPUT3), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n376), .A2(new_n331), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n434), .C1(new_n436), .C2(new_n344), .ZN(new_n437));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n365), .B1(new_n430), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n394), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n351), .B2(new_n435), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n437), .A2(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT82), .B(G22gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  XOR2_X1   g248(.A(new_n449), .B(KEYINPUT79), .Z(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n444), .B2(new_n445), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n446), .A2(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n364), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n353), .A2(new_n358), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n345), .A2(new_n352), .A3(KEYINPUT30), .A4(new_n363), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n401), .A2(new_n392), .A3(new_n402), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT39), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(KEYINPUT84), .A3(KEYINPUT39), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n406), .A2(new_n391), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n392), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n392), .B1(new_n406), .B2(new_n391), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n415), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n461), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n416), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n473), .B2(new_n472), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n454), .B1(new_n460), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n429), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n397), .B(new_n292), .C1(new_n328), .C2(new_n329), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n321), .A2(new_n312), .A3(new_n308), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT70), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n397), .A4(new_n292), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n330), .A2(new_n395), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n485), .B(KEYINPUT64), .Z(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT65), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n484), .A2(KEYINPUT34), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT34), .B1(new_n484), .B2(new_n486), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n484), .A2(new_n487), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT71), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n487), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G71gat), .B(G99gat), .Z(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G43gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT33), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n490), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n487), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT71), .B1(new_n484), .B2(new_n487), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT32), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT33), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n506), .A3(new_n499), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n496), .A2(new_n500), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n507), .A2(new_n509), .B1(new_n489), .B2(new_n488), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT36), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n508), .A2(new_n510), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT78), .A4(new_n412), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n405), .A2(new_n407), .A3(new_n412), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n414), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n418), .ZN(new_n520));
  AND4_X1   g319(.A1(new_n520), .A2(new_n456), .A3(new_n459), .A4(new_n457), .ZN(new_n521));
  INV_X1    g320(.A(new_n454), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n477), .A2(new_n511), .A3(new_n514), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n490), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n454), .B1(new_n501), .B2(new_n507), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT35), .B1(new_n417), .B2(new_n418), .ZN(new_n530));
  AND4_X1   g329(.A1(new_n459), .A2(new_n530), .A3(new_n457), .A4(new_n456), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n526), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n271), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G64gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(G57gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(G57gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(KEYINPUT98), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(KEYINPUT98), .B2(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  OR2_X1    g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n537), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT9), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n540), .A3(new_n541), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n549));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(G127gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n259), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n553), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT99), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G155gat), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n556), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n576), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n572), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT100), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n251), .A2(new_n252), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n577), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n582), .A2(new_n242), .B1(KEYINPUT41), .B2(new_n564), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT101), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n586), .A3(new_n583), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n585), .B2(new_n587), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n568), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n567), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n548), .B1(new_n580), .B2(new_n577), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n544), .A2(new_n547), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n579), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n602), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n582), .A2(KEYINPUT10), .A3(new_n548), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n603), .A2(new_n605), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n601), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(KEYINPUT102), .A3(new_n600), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND4_X1   g419(.A1(new_n534), .A2(new_n563), .A3(new_n597), .A4(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n520), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G1gat), .ZN(G1324gat));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n460), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT103), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT16), .B(G8gat), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(G8gat), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n626), .A2(new_n625), .A3(new_n628), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(G1325gat));
  AOI21_X1  g431(.A(G15gat), .B1(new_n621), .B2(new_n512), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n514), .A2(new_n511), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(G15gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT104), .Z(new_n636));
  AOI21_X1  g435(.A(new_n633), .B1(new_n621), .B2(new_n636), .ZN(G1326gat));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n454), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT43), .B(G22gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1327gat));
  AND2_X1   g439(.A1(new_n524), .A2(new_n533), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n562), .A2(new_n620), .ZN(new_n642));
  NOR4_X1   g441(.A1(new_n641), .A2(new_n271), .A3(new_n597), .A4(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G29gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n622), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT105), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT45), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n529), .A2(KEYINPUT106), .A3(new_n532), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT106), .B1(new_n529), .B2(new_n532), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n524), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n524), .B(KEYINPUT107), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n597), .A2(KEYINPUT44), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT44), .B1(new_n641), .B2(new_n597), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n271), .B(new_n642), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n659), .A2(new_n622), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n648), .B(new_n649), .C1(new_n644), .C2(new_n660), .ZN(G1328gat));
  INV_X1    g460(.A(G36gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n643), .A2(new_n662), .A3(new_n460), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(KEYINPUT108), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(KEYINPUT108), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n659), .A2(new_n460), .ZN(new_n668));
  OAI221_X1 g467(.A(new_n667), .B1(new_n665), .B2(new_n663), .C1(new_n668), .C2(new_n662), .ZN(G1329gat));
  NAND2_X1  g468(.A1(new_n659), .A2(new_n634), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n508), .A2(new_n510), .A3(G43gat), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n670), .A2(G43gat), .B1(new_n643), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n643), .B2(new_n454), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n454), .A2(G50gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n659), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1331gat));
  AND2_X1   g477(.A1(new_n654), .A2(new_n655), .ZN(new_n679));
  NOR4_X1   g478(.A1(new_n596), .A2(new_n270), .A3(new_n562), .A4(new_n620), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n622), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G57gat), .ZN(G1332gat));
  INV_X1    g482(.A(new_n460), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT110), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n687), .B(KEYINPUT111), .ZN(new_n692));
  INV_X1    g491(.A(new_n690), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(G1333gat));
  NAND2_X1  g494(.A1(new_n681), .A2(new_n634), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G71gat), .ZN(new_n697));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n698), .A3(new_n512), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1334gat));
  NAND2_X1  g501(.A1(new_n681), .A2(new_n454), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g503(.A1(new_n270), .A2(new_n563), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n619), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n657), .B2(new_n658), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G85gat), .B1(new_n708), .B2(new_n520), .ZN(new_n709));
  INV_X1    g508(.A(new_n705), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n533), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n529), .A2(KEYINPUT106), .A3(new_n532), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n597), .B1(new_n714), .B2(new_n524), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n710), .B1(new_n715), .B2(KEYINPUT113), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT113), .B1(new_n652), .B2(new_n596), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT51), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n652), .A2(KEYINPUT113), .A3(new_n596), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n705), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n619), .A2(new_n574), .A3(new_n622), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n709), .B1(new_n724), .B2(new_n725), .ZN(G1336gat));
  AOI21_X1  g525(.A(new_n575), .B1(new_n707), .B2(new_n460), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT52), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n460), .A2(new_n575), .A3(new_n619), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n722), .B2(new_n717), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n729), .B1(new_n719), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT52), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(G1337gat));
  INV_X1    g535(.A(new_n634), .ZN(new_n737));
  OAI21_X1  g536(.A(G99gat), .B1(new_n708), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(G99gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n512), .A2(new_n739), .A3(new_n619), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n724), .B2(new_n740), .ZN(G1338gat));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n620), .A2(G106gat), .A3(new_n522), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n719), .B2(new_n723), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT115), .B(G106gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n707), .B2(new_n454), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT53), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n731), .B1(new_n716), .B2(new_n718), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n722), .A2(new_n720), .A3(new_n717), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n657), .A2(new_n658), .ZN(new_n753));
  INV_X1    g552(.A(new_n706), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n454), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n746), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n742), .B1(new_n748), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n744), .B1(new_n719), .B2(new_n733), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT53), .B1(new_n760), .B2(new_n747), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n749), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n761), .B(KEYINPUT116), .C1(new_n745), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(G1339gat));
  NOR4_X1   g563(.A1(new_n596), .A2(new_n270), .A3(new_n562), .A4(new_n619), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n601), .B1(new_n610), .B2(KEYINPUT54), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT118), .B(new_n601), .C1(new_n610), .C2(KEYINPUT54), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n606), .A2(new_n612), .A3(new_n607), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n610), .A2(KEYINPUT54), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT117), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n610), .A2(new_n774), .A3(KEYINPUT54), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n615), .A2(new_n600), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n770), .A2(KEYINPUT55), .A3(new_n776), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n262), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n248), .A2(new_n260), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n249), .B1(new_n248), .B2(new_n253), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n205), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n256), .A2(new_n263), .A3(new_n207), .A4(new_n258), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n596), .A2(new_n782), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n787), .A2(new_n619), .A3(new_n786), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n270), .B2(new_n782), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(new_n596), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n765), .B1(new_n791), .B2(new_n562), .ZN(new_n792));
  NOR4_X1   g591(.A1(new_n792), .A2(new_n510), .A3(new_n508), .A4(new_n454), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n622), .A3(new_n684), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n271), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n620), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g597(.A1(new_n794), .A2(new_n562), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n552), .A2(KEYINPUT119), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n799), .B(new_n800), .Z(G1342gat));
  NOR2_X1   g600(.A1(new_n597), .A2(new_n460), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n520), .A2(G134gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n793), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT56), .Z(new_n805));
  OAI21_X1  g604(.A(G134gat), .B1(new_n794), .B2(new_n597), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1343gat));
  OAI21_X1  g606(.A(KEYINPUT57), .B1(new_n792), .B2(new_n522), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n269), .B2(new_n265), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n597), .B1(new_n811), .B2(new_n789), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n563), .B1(new_n812), .B2(new_n788), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n809), .B(new_n454), .C1(new_n813), .C2(new_n765), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n634), .A2(new_n520), .A3(new_n460), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n808), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G141gat), .B1(new_n816), .B2(new_n271), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818));
  INV_X1    g617(.A(new_n792), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n454), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n634), .A2(new_n520), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n684), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n271), .A2(G141gat), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n817), .B(new_n818), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n816), .A2(KEYINPUT120), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n808), .A2(new_n814), .A3(new_n829), .A4(new_n815), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n270), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n824), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n831), .A2(G141gat), .B1(new_n832), .B2(new_n825), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n833), .B2(new_n818), .ZN(G1344gat));
  NAND3_X1  g633(.A1(new_n828), .A2(new_n619), .A3(new_n830), .ZN(new_n835));
  INV_X1    g634(.A(G148gat), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT59), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n808), .A2(new_n814), .A3(new_n619), .A4(new_n815), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G148gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT59), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n838), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n619), .A2(new_n836), .ZN(new_n846));
  OR3_X1    g645(.A1(new_n824), .A2(KEYINPUT121), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT121), .B1(new_n824), .B2(new_n846), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(G1345gat));
  AOI21_X1  g649(.A(G155gat), .B1(new_n832), .B2(new_n563), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n828), .A2(new_n830), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n563), .A2(G155gat), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT123), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(G1346gat));
  INV_X1    g654(.A(G162gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n823), .A2(new_n856), .A3(new_n802), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n852), .A2(new_n596), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n856), .ZN(G1347gat));
  NOR2_X1   g658(.A1(new_n684), .A2(new_n622), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n793), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n271), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT124), .B(G169gat), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(G1348gat));
  NOR2_X1   g663(.A1(new_n861), .A2(new_n620), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT125), .B(G176gat), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(G1349gat));
  OAI21_X1  g666(.A(new_n303), .B1(new_n861), .B2(new_n562), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n793), .A2(new_n286), .A3(new_n563), .A4(new_n860), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(G1350gat));
  OAI22_X1  g671(.A1(new_n861), .A2(new_n597), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n873), .B(new_n874), .ZN(G1351gat));
  AND2_X1   g674(.A1(new_n808), .A2(new_n814), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n634), .A2(new_n622), .A3(new_n684), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(G197gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n878), .A2(new_n879), .A3(new_n271), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n819), .A2(new_n454), .A3(new_n877), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(new_n271), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n879), .B2(new_n882), .ZN(G1352gat));
  OAI21_X1  g682(.A(G204gat), .B1(new_n878), .B2(new_n620), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n620), .A2(G204gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886));
  OAI22_X1  g685(.A1(new_n881), .A2(new_n885), .B1(new_n886), .B2(KEYINPUT62), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(KEYINPUT126), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n886), .B(KEYINPUT62), .C1(new_n881), .C2(new_n885), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(G1353gat));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n563), .A3(new_n877), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n336), .B1(KEYINPUT127), .B2(new_n895), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n893), .A2(new_n896), .B1(new_n892), .B2(KEYINPUT63), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n563), .A2(new_n336), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n894), .A2(new_n897), .B1(new_n881), .B2(new_n898), .ZN(G1354gat));
  OAI21_X1  g698(.A(G218gat), .B1(new_n878), .B2(new_n597), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n596), .A2(new_n337), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n881), .B2(new_n901), .ZN(G1355gat));
endmodule


