//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n458), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G124), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n458), .A2(G112), .ZN(new_n473));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n471), .A2(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n458), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(KEYINPUT65), .A3(new_n458), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n475), .B1(new_n480), .B2(G136), .ZN(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(KEYINPUT66), .B2(G114), .ZN(new_n483));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G114), .ZN(new_n484));
  OAI211_X1 g059(.A(G2104), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n460), .A2(new_n462), .A3(G126), .A4(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT67), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n458), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n470), .A2(new_n493), .A3(G138), .A4(new_n458), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n488), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT68), .A3(G50), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n499), .A2(new_n501), .A3(new_n511), .A4(new_n513), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n515), .A2(new_n498), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n509), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT69), .B(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n503), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n520), .B(KEYINPUT70), .C1(new_n503), .C2(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  INV_X1    g103(.A(new_n517), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n528), .B1(new_n529), .B2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n511), .A2(new_n513), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n529), .A2(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n503), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n504), .A2(G52), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n543), .A2(KEYINPUT71), .A3(new_n537), .A4(new_n538), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n534), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n503), .A2(new_n551), .B1(new_n552), .B2(new_n517), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n502), .A2(new_n514), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G91), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n499), .A2(new_n501), .A3(G53), .A4(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n534), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n568), .A2(new_n569), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n566), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n526), .A2(new_n577), .A3(new_n530), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND2_X1  g155(.A1(new_n565), .A2(G87), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n498), .B1(new_n534), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n504), .B2(G49), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT74), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT74), .B1(new_n581), .B2(new_n584), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT75), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n511), .A2(new_n513), .A3(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n498), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(G48), .A2(new_n504), .B1(new_n594), .B2(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n565), .A2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n593), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n498), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n503), .A2(new_n604), .B1(new_n605), .B2(new_n517), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n565), .A2(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n534), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n504), .A2(G54), .B1(new_n615), .B2(G651), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n609), .B1(new_n618), .B2(G868), .ZN(G321));
  XNOR2_X1  g194(.A(G321), .B(KEYINPUT77), .ZN(G284));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(G868), .B2(new_n622), .ZN(G297));
  OAI21_X1  g198(.A(new_n621), .B1(G868), .B2(new_n622), .ZN(G280));
  INV_X1    g199(.A(G860), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n617), .B1(G559), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT78), .ZN(G148));
  OR2_X1    g202(.A1(new_n617), .A2(G559), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(new_n471), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G123), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n480), .B2(G135), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT79), .B(G2096), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n458), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT16), .B(G1341), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(G14), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n651), .A2(new_n657), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(KEYINPUT81), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n662), .B(KEYINPUT17), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n667), .B2(new_n663), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(KEYINPUT81), .B2(new_n664), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  INV_X1    g245(.A(new_n661), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n671), .A2(new_n662), .A3(new_n663), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n667), .A2(new_n661), .A3(new_n663), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n685), .B1(new_n683), .B2(new_n681), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1991), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT85), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(G229));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT26), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n458), .A2(G105), .A3(G2104), .ZN(new_n702));
  INV_X1    g277(.A(G129), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n701), .B(new_n702), .C1(new_n471), .C2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G141), .B2(new_n480), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT97), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G29), .B2(G32), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G33), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT25), .Z(new_n714));
  AOI22_X1  g289(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n458), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n480), .B2(G139), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(new_n711), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2072), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G5), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G171), .B2(new_n720), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G1961), .ZN(new_n723));
  NOR2_X1   g298(.A1(G164), .A2(new_n711), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G27), .B2(new_n711), .ZN(new_n725));
  INV_X1    g300(.A(G2078), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n722), .A2(G1961), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n719), .A2(new_n723), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1956), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n720), .A2(G20), .ZN(new_n731));
  NAND2_X1  g306(.A1(G299), .A2(G16), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(KEYINPUT23), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(KEYINPUT23), .B2(new_n731), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n710), .B(new_n735), .C1(new_n730), .C2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT28), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n711), .A2(G26), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n480), .A2(G140), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n480), .A2(KEYINPUT94), .A3(G140), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G116), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n632), .A2(G128), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n741), .A2(new_n742), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n737), .B(new_n738), .C1(new_n748), .C2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n737), .B2(new_n738), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT96), .B(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n618), .B2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT91), .B(G1348), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n555), .A2(new_n720), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n720), .B2(G19), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT92), .B(G1341), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G160), .B2(new_n711), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n759), .A2(new_n761), .B1(G2084), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G2084), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n637), .A2(G29), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G28), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n711), .B1(new_n770), .B2(G28), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AND2_X1   g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n769), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n759), .B2(new_n761), .ZN(new_n776));
  NAND2_X1  g351(.A1(G168), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G16), .B2(G21), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(new_n726), .B2(new_n725), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n757), .A2(new_n768), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n778), .A2(new_n779), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT98), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2090), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n711), .A2(G35), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G162), .B2(new_n711), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT29), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n784), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(G2090), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n782), .A2(new_n783), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n781), .A2(new_n790), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n736), .A2(new_n752), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n720), .A2(G6), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n499), .A2(new_n501), .A3(G48), .A4(G543), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n598), .B2(new_n599), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n594), .A2(KEYINPUT76), .ZN(new_n799));
  INV_X1    g374(.A(G86), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n563), .B2(new_n564), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n720), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n720), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n720), .ZN(new_n810));
  INV_X1    g385(.A(G1971), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G23), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n581), .A2(new_n584), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT33), .B(G1976), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n807), .A2(new_n808), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT34), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n711), .A2(G25), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n632), .A2(KEYINPUT86), .A3(G119), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT86), .ZN(new_n822));
  INV_X1    g397(.A(G119), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n471), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g399(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT87), .B1(G95), .B2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n821), .B(new_n824), .C1(new_n825), .C2(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n480), .A2(G131), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n820), .B1(new_n830), .B2(new_n711), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n720), .A2(G24), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n607), .B2(new_n720), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1986), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n819), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT90), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(KEYINPUT90), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n838), .A2(KEYINPUT90), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n795), .B1(new_n843), .B2(new_n844), .ZN(G311));
  INV_X1    g420(.A(new_n795), .ZN(new_n846));
  INV_X1    g421(.A(new_n842), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n841), .B1(new_n838), .B2(KEYINPUT90), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(new_n618), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n852));
  XOR2_X1   g427(.A(new_n851), .B(new_n852), .Z(new_n853));
  AOI22_X1  g428(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n498), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n503), .A2(new_n856), .B1(new_n857), .B2(new_n517), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n554), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n853), .A2(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n625), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(G162), .B(KEYINPUT100), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G160), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n637), .B(new_n705), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n748), .B(new_n641), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT101), .B1(new_n458), .B2(G118), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n458), .A2(KEYINPUT101), .A3(G118), .ZN(new_n875));
  INV_X1    g450(.A(G130), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n874), .A2(new_n875), .B1(new_n471), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n480), .B2(G142), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n485), .A2(new_n486), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n495), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n878), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n872), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n871), .B(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n830), .B(new_n717), .Z(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g464(.A(new_n628), .B(new_n861), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n617), .A2(new_n622), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n612), .A2(G299), .A3(new_n616), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n895), .B1(new_n890), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G305), .B(new_n607), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(G303), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n814), .B(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(G303), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n905), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n901), .A2(new_n902), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n903), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n903), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n859), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(G868), .B2(new_n915), .ZN(G295));
  OAI21_X1  g491(.A(new_n914), .B1(G868), .B2(new_n915), .ZN(G331));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(G301), .A2(new_n531), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n861), .B(new_n920), .C1(G286), .C2(G301), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(new_n894), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(G286), .B2(G301), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n924), .A2(new_n860), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n860), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n923), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n921), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n931), .A2(new_n900), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n931), .B2(new_n900), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n930), .B(new_n910), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n886), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n894), .A2(new_n896), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n893), .A2(new_n898), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n927), .B(KEYINPUT105), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n922), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n923), .A2(new_n927), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n910), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n919), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n910), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n938), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n927), .B(new_n928), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(new_n921), .ZN(new_n947));
  INV_X1    g522(.A(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n949), .A2(KEYINPUT106), .A3(new_n886), .A4(new_n935), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n918), .B1(new_n943), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n936), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n944), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n918), .B1(new_n952), .B2(new_n954), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n936), .A2(new_n942), .A3(KEYINPUT43), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(G397));
  INV_X1    g536(.A(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n495), .B2(new_n879), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(KEYINPUT107), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G160), .A2(G40), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n705), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(G1996), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n974));
  INV_X1    g549(.A(G2067), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n748), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G1996), .B2(new_n971), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n973), .B(new_n974), .C1(new_n977), .C2(new_n970), .ZN(new_n978));
  INV_X1    g553(.A(new_n970), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n830), .B(new_n832), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT108), .ZN(new_n983));
  NAND2_X1  g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  AOI22_X1  g563(.A1(KEYINPUT67), .A2(new_n487), .B1(new_n492), .B2(new_n494), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n989), .B2(new_n490), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n496), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n969), .B1(new_n963), .B2(new_n991), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n992), .A2(new_n785), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n969), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n811), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G8), .B1(new_n509), .B2(new_n518), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(G8), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1003), .A2(KEYINPUT111), .A3(G8), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n465), .A2(new_n468), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n963), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n814), .B2(G1976), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n585), .B2(new_n586), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n797), .B1(new_n517), .B2(new_n800), .ZN(new_n1022));
  OAI21_X1  g597(.A(G1981), .B1(new_n1022), .B2(new_n594), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT112), .B(G1981), .C1(new_n1022), .C2(new_n594), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n595), .A2(new_n596), .A3(new_n1028), .A4(new_n600), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1015), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT49), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1030), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT114), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n1037), .B2(KEYINPUT49), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1021), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1002), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n496), .A2(new_n991), .A3(new_n993), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1013), .B1(new_n963), .B2(new_n991), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1045), .A2(new_n1046), .A3(G2090), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1006), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G2084), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n992), .A2(new_n1051), .A3(new_n995), .A4(new_n996), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n994), .A2(new_n998), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1013), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n779), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G286), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1011), .A2(new_n1043), .A3(new_n1050), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1006), .B1(new_n1003), .B2(G8), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1062), .A2(new_n1057), .A3(new_n1060), .A4(G286), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(new_n1011), .A3(new_n1043), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1066));
  OR2_X1    g641(.A1(G288), .A2(G1976), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1029), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1011), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1068), .A2(new_n1031), .B1(new_n1069), .B2(new_n1043), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(G8), .C1(new_n1056), .C2(new_n531), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n531), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT123), .B1(new_n1056), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1077), .B(new_n1074), .C1(new_n1052), .C2(new_n1055), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1073), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1072), .B(new_n1075), .C1(new_n1056), .C2(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1056), .A2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1077), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1056), .A2(KEYINPUT123), .A3(new_n1075), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1057), .A2(KEYINPUT51), .A3(new_n1074), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1073), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1054), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n726), .C1(new_n998), .C2(new_n994), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n1095));
  INV_X1    g670(.A(G1961), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n999), .A2(new_n726), .A3(new_n1000), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1095), .A2(new_n1096), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1081), .A2(new_n1088), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1011), .A2(new_n1043), .A3(new_n1050), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1011), .A2(new_n1043), .A3(KEYINPUT126), .A4(new_n1050), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1071), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n991), .B1(new_n496), .B2(new_n993), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n996), .B1(new_n1107), .B2(KEYINPUT110), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n990), .A2(new_n988), .A3(new_n991), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n756), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1014), .B2(G2067), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n963), .A2(new_n1013), .A3(KEYINPUT118), .A4(new_n975), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n1115), .A4(new_n617), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n618), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1114), .B1(new_n1095), .B2(new_n756), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n617), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1120), .A2(KEYINPUT60), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1001), .A2(G1996), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n963), .B2(new_n1013), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n555), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT59), .B(new_n555), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT115), .B(G1956), .Z(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(G2072), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n999), .A2(new_n1000), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n568), .B2(new_n569), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G299), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n566), .B(new_n573), .C1(new_n1140), .C2(KEYINPUT57), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1135), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1132), .B(new_n1133), .C1(new_n1148), .C2(KEYINPUT61), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1147), .B2(KEYINPUT119), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1135), .A2(new_n1138), .A3(new_n1144), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(KEYINPUT61), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1150), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1152), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1123), .A2(new_n1158), .A3(new_n1124), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1126), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1120), .A2(new_n617), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1145), .B1(new_n1161), .B2(new_n1147), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1164));
  XOR2_X1   g739(.A(G171), .B(KEYINPUT54), .Z(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT53), .B1(new_n1166), .B2(G2078), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1166), .B2(G2078), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1000), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1165), .B1(new_n968), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1164), .A2(new_n1165), .B1(new_n1170), .B2(new_n1098), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n987), .B1(new_n1106), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n979), .A2(new_n983), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT48), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n981), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  OR3_X1    g754(.A1(new_n979), .A2(new_n1179), .A3(G1996), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n979), .B2(G1996), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n976), .A2(new_n705), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1180), .B(new_n1181), .C1(new_n1182), .C2(new_n979), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n828), .A2(new_n829), .A3(new_n832), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n978), .A2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n748), .A2(G2067), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1178), .B(new_n1184), .C1(new_n979), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n962), .B1(new_n1175), .B2(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1065), .B(new_n1070), .C1(new_n1192), .C2(new_n1100), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n986), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1188), .A2(new_n979), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1194), .A2(new_n1197), .A3(KEYINPUT127), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1190), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g774(.A1(new_n958), .A2(new_n959), .ZN(new_n1201));
  OAI21_X1  g775(.A(G319), .B1(new_n658), .B2(new_n659), .ZN(new_n1202));
  NOR3_X1   g776(.A1(G229), .A2(G227), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g777(.A(new_n1203), .B1(new_n887), .B2(new_n885), .ZN(new_n1204));
  NOR2_X1   g778(.A1(new_n1201), .A2(new_n1204), .ZN(G308));
  INV_X1    g779(.A(G308), .ZN(G225));
endmodule


