

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n463), .B(n462), .ZN(n523) );
  AND2_X1 U322 ( .A1(G227GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n454) );
  XNOR2_X1 U324 ( .A(n455), .B(n454), .ZN(n461) );
  XNOR2_X1 U325 ( .A(n523), .B(KEYINPUT115), .ZN(n464) );
  INV_X1 U326 ( .A(KEYINPUT48), .ZN(n462) );
  XNOR2_X1 U327 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U328 ( .A(n298), .B(n289), .ZN(n299) );
  XNOR2_X1 U329 ( .A(n424), .B(n423), .ZN(n428) );
  XNOR2_X1 U330 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n407) );
  XNOR2_X1 U331 ( .A(n371), .B(n299), .ZN(n307) );
  XNOR2_X1 U332 ( .A(n408), .B(n407), .ZN(n512) );
  NOR2_X1 U333 ( .A1(n528), .A2(n469), .ZN(n561) );
  INV_X1 U334 ( .A(G43GAT), .ZN(n447) );
  XNOR2_X1 U335 ( .A(n396), .B(n308), .ZN(n528) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n470) );
  XNOR2_X1 U337 ( .A(n447), .B(KEYINPUT40), .ZN(n448) );
  XNOR2_X1 U338 ( .A(n471), .B(n470), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n449), .B(n448), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT0), .B(KEYINPUT78), .Z(n291) );
  XNOR2_X1 U341 ( .A(KEYINPUT77), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U343 ( .A(G113GAT), .B(n292), .Z(n396) );
  XOR2_X1 U344 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U345 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U347 ( .A(G169GAT), .B(n295), .Z(n371) );
  XOR2_X1 U348 ( .A(G134GAT), .B(G190GAT), .Z(n297) );
  XNOR2_X1 U349 ( .A(KEYINPUT79), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U351 ( .A(KEYINPUT20), .B(G71GAT), .Z(n301) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G176GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U354 ( .A(G183GAT), .B(KEYINPUT80), .Z(n303) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G99GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(n305), .B(n304), .Z(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U359 ( .A(G71GAT), .B(KEYINPUT13), .Z(n420) );
  XOR2_X1 U360 ( .A(G1GAT), .B(KEYINPUT67), .Z(n310) );
  XNOR2_X1 U361 ( .A(G22GAT), .B(G15GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n431) );
  XOR2_X1 U363 ( .A(n420), .B(n431), .Z(n312) );
  NAND2_X1 U364 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(n313), .B(KEYINPUT15), .Z(n316) );
  XNOR2_X1 U367 ( .A(G8GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n314), .B(KEYINPUT74), .ZN(n369) );
  XNOR2_X1 U369 ( .A(G57GAT), .B(n369), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n324) );
  XOR2_X1 U371 ( .A(G78GAT), .B(G155GAT), .Z(n318) );
  XNOR2_X1 U372 ( .A(G127GAT), .B(G211GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U374 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n320) );
  XNOR2_X1 U375 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U377 ( .A(n322), .B(n321), .Z(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n578) );
  INV_X1 U379 ( .A(n578), .ZN(n456) );
  XNOR2_X1 U380 ( .A(G218GAT), .B(G106GAT), .ZN(n325) );
  XOR2_X1 U381 ( .A(G36GAT), .B(G190GAT), .Z(n364) );
  XNOR2_X1 U382 ( .A(n325), .B(n364), .ZN(n339) );
  XNOR2_X1 U383 ( .A(G29GAT), .B(G134GAT), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n326), .B(KEYINPUT73), .ZN(n381) );
  XOR2_X1 U385 ( .A(G92GAT), .B(n381), .Z(n328) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U388 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n330) );
  XNOR2_X1 U389 ( .A(G162GAT), .B(KEYINPUT10), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U391 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U392 ( .A(G43GAT), .B(G50GAT), .Z(n334) );
  XNOR2_X1 U393 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n442) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G85GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n335), .B(KEYINPUT70), .ZN(n425) );
  XNOR2_X1 U397 ( .A(n442), .B(n425), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n552) );
  INV_X1 U400 ( .A(n552), .ZN(n473) );
  XNOR2_X1 U401 ( .A(KEYINPUT36), .B(n473), .ZN(n580) );
  XOR2_X1 U402 ( .A(KEYINPUT84), .B(G218GAT), .Z(n341) );
  XNOR2_X1 U403 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U405 ( .A(G197GAT), .B(n342), .Z(n370) );
  XOR2_X1 U406 ( .A(G148GAT), .B(KEYINPUT83), .Z(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT82), .B(KEYINPUT23), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U409 ( .A(G106GAT), .B(G78GAT), .Z(n409) );
  XOR2_X1 U410 ( .A(n345), .B(n409), .Z(n347) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G22GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U413 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n349) );
  NAND2_X1 U414 ( .A1(G228GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U416 ( .A(n351), .B(n350), .Z(n357) );
  XNOR2_X1 U417 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n352), .B(KEYINPUT2), .ZN(n353) );
  XOR2_X1 U419 ( .A(n353), .B(KEYINPUT85), .Z(n355) );
  XNOR2_X1 U420 ( .A(G141GAT), .B(G162GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n391) );
  XNOR2_X1 U422 ( .A(n391), .B(G204GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n370), .B(n358), .ZN(n467) );
  NAND2_X1 U425 ( .A1(n467), .A2(n528), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n359), .B(KEYINPUT94), .ZN(n360) );
  XNOR2_X1 U427 ( .A(KEYINPUT26), .B(n360), .ZN(n563) );
  XOR2_X1 U428 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n362) );
  XNOR2_X1 U429 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U431 ( .A(n364), .B(n363), .Z(n366) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n375) );
  XOR2_X1 U434 ( .A(G64GAT), .B(G92GAT), .Z(n368) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G204GAT), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n368), .B(n367), .ZN(n426) );
  XOR2_X1 U437 ( .A(n369), .B(n426), .Z(n373) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U440 ( .A(n375), .B(n374), .Z(n516) );
  XNOR2_X1 U441 ( .A(n516), .B(KEYINPUT27), .ZN(n402) );
  NOR2_X1 U442 ( .A1(n563), .A2(n402), .ZN(n380) );
  NOR2_X1 U443 ( .A1(n528), .A2(n516), .ZN(n376) );
  NOR2_X1 U444 ( .A1(n467), .A2(n376), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n377), .B(KEYINPUT25), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n378), .B(KEYINPUT95), .ZN(n379) );
  NOR2_X1 U447 ( .A1(n380), .A2(n379), .ZN(n399) );
  XOR2_X1 U448 ( .A(n381), .B(KEYINPUT1), .Z(n383) );
  NAND2_X1 U449 ( .A1(G225GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U454 ( .A(G85GAT), .B(KEYINPUT6), .Z(n387) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(KEYINPUT87), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U457 ( .A(n389), .B(n388), .Z(n393) );
  XNOR2_X1 U458 ( .A(G120GAT), .B(G148GAT), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n390), .B(G57GAT), .ZN(n410) );
  XNOR2_X1 U460 ( .A(n391), .B(n410), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n398) );
  INV_X1 U463 ( .A(n396), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n401) );
  NOR2_X1 U465 ( .A1(n399), .A2(n401), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT96), .ZN(n405) );
  XNOR2_X1 U467 ( .A(KEYINPUT89), .B(n401), .ZN(n565) );
  NOR2_X1 U468 ( .A1(n565), .A2(n402), .ZN(n524) );
  NAND2_X1 U469 ( .A1(n528), .A2(n524), .ZN(n403) );
  XNOR2_X1 U470 ( .A(KEYINPUT28), .B(n467), .ZN(n526) );
  NOR2_X1 U471 ( .A1(n403), .A2(n526), .ZN(n404) );
  NOR2_X1 U472 ( .A1(n405), .A2(n404), .ZN(n477) );
  NOR2_X1 U473 ( .A1(n580), .A2(n477), .ZN(n406) );
  NAND2_X1 U474 ( .A1(n456), .A2(n406), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  AND2_X1 U476 ( .A1(G230GAT), .A2(G233GAT), .ZN(n412) );
  NAND2_X1 U477 ( .A1(n411), .A2(n412), .ZN(n416) );
  INV_X1 U478 ( .A(n411), .ZN(n414) );
  INV_X1 U479 ( .A(n412), .ZN(n413) );
  NAND2_X1 U480 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U481 ( .A1(n416), .A2(n415), .ZN(n417) );
  XOR2_X1 U482 ( .A(n417), .B(KEYINPUT69), .Z(n424) );
  XOR2_X1 U483 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n419) );
  XNOR2_X1 U484 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n418) );
  XOR2_X1 U485 ( .A(n419), .B(n418), .Z(n422) );
  XNOR2_X1 U486 ( .A(n420), .B(KEYINPUT32), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n573) );
  XOR2_X1 U489 ( .A(G36GAT), .B(G29GAT), .Z(n430) );
  NAND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U492 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U493 ( .A(G113GAT), .B(G141GAT), .Z(n434) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(G197GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n436) );
  XNOR2_X1 U497 ( .A(G8GAT), .B(KEYINPUT66), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U501 ( .A(n441), .B(KEYINPUT65), .Z(n444) );
  XNOR2_X1 U502 ( .A(n442), .B(KEYINPUT64), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n569) );
  NAND2_X1 U504 ( .A1(n573), .A2(n569), .ZN(n445) );
  XOR2_X1 U505 ( .A(KEYINPUT72), .B(n445), .Z(n479) );
  NAND2_X1 U506 ( .A1(n512), .A2(n479), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n446), .B(KEYINPUT38), .ZN(n498) );
  NOR2_X1 U508 ( .A1(n528), .A2(n498), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n573), .B(KEYINPUT41), .ZN(n544) );
  NAND2_X1 U510 ( .A1(n544), .A2(n569), .ZN(n451) );
  XOR2_X1 U511 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n450) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(n453) );
  NOR2_X1 U513 ( .A1(n552), .A2(n578), .ZN(n452) );
  NAND2_X1 U514 ( .A1(n453), .A2(n452), .ZN(n455) );
  NOR2_X1 U515 ( .A1(n456), .A2(n580), .ZN(n457) );
  XNOR2_X1 U516 ( .A(KEYINPUT45), .B(n457), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n458), .A2(n573), .ZN(n459) );
  NOR2_X1 U518 ( .A1(n459), .A2(n569), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n464), .A2(n516), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT54), .ZN(n567) );
  NAND2_X1 U522 ( .A1(n567), .A2(n565), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT55), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n552), .A2(n561), .ZN(n471) );
  XOR2_X1 U526 ( .A(G1GAT), .B(KEYINPUT34), .Z(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT99), .B(n472), .ZN(n482) );
  NAND2_X1 U528 ( .A1(n578), .A2(n473), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT76), .ZN(n475) );
  XNOR2_X1 U530 ( .A(n475), .B(KEYINPUT16), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U532 ( .A(KEYINPUT97), .B(n478), .Z(n501) );
  NAND2_X1 U533 ( .A1(n479), .A2(n501), .ZN(n480) );
  XNOR2_X1 U534 ( .A(n480), .B(KEYINPUT98), .ZN(n487) );
  NOR2_X1 U535 ( .A1(n565), .A2(n487), .ZN(n481) );
  XOR2_X1 U536 ( .A(n482), .B(n481), .Z(G1324GAT) );
  NOR2_X1 U537 ( .A1(n516), .A2(n487), .ZN(n483) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n485) );
  NOR2_X1 U540 ( .A1(n528), .A2(n487), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n526), .ZN(n520) );
  NOR2_X1 U544 ( .A1(n487), .A2(n520), .ZN(n489) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n492) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n494) );
  NOR2_X1 U551 ( .A1(n565), .A2(n498), .ZN(n493) );
  XOR2_X1 U552 ( .A(n494), .B(n493), .Z(G1328GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n496) );
  NOR2_X1 U554 ( .A1(n516), .A2(n498), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U557 ( .A1(n498), .A2(n520), .ZN(n499) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  XNOR2_X1 U559 ( .A(KEYINPUT108), .B(n544), .ZN(n558) );
  INV_X1 U560 ( .A(n558), .ZN(n500) );
  NOR2_X1 U561 ( .A1(n569), .A2(n500), .ZN(n513) );
  NAND2_X1 U562 ( .A1(n501), .A2(n513), .ZN(n508) );
  NOR2_X1 U563 ( .A1(n565), .A2(n508), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(n502), .Z(n503) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n516), .A2(n508), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n528), .A2(n508), .ZN(n506) );
  XOR2_X1 U570 ( .A(KEYINPUT110), .B(n506), .Z(n507) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U572 ( .A1(n520), .A2(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U575 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n519) );
  NOR2_X1 U577 ( .A1(n565), .A2(n519), .ZN(n514) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT112), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n519), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n530) );
  XOR2_X1 U588 ( .A(KEYINPUT115), .B(n523), .Z(n525) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n539) );
  OR2_X1 U590 ( .A1(n539), .A2(n526), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n569), .A2(n536), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U595 ( .A1(n536), .A2(n558), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NAND2_X1 U598 ( .A1(n578), .A2(n536), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U602 ( .A1(n536), .A2(n552), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U604 ( .A1(n563), .A2(n539), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n569), .A2(n551), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT118), .B(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n543) );
  XNOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n548) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n578), .A2(n551), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT122), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n561), .A2(n569), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(n557), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n578), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  INV_X1 U631 ( .A(n563), .ZN(n564) );
  AND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(n568), .Z(n577) );
  NAND2_X1 U635 ( .A1(n577), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  INV_X1 U638 ( .A(n577), .ZN(n581) );
  OR2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

