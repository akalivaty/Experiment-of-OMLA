//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n188), .B(G101), .ZN(new_n193));
  INV_X1    g007(.A(new_n191), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n192), .A2(new_n195), .A3(KEYINPUT67), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT67), .B1(new_n192), .B2(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT2), .A2(G113), .ZN(new_n206));
  XNOR2_X1  g020(.A(G116), .B(G119), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT0), .B(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G137), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n222), .A2(new_n224), .A3(new_n228), .A4(new_n225), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n219), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n213), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n211), .A2(G143), .ZN(new_n233));
  OAI211_X1 g047(.A(G128), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n221), .A2(G137), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n223), .A2(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(G131), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n212), .B(new_n214), .C1(KEYINPUT1), .C2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n234), .A2(new_n229), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n210), .B1(new_n230), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n227), .A2(new_n229), .ZN(new_n243));
  INV_X1    g057(.A(new_n219), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n208), .A2(new_n209), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n240), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n199), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n247), .A2(new_n199), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n198), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n192), .A2(new_n195), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n230), .B2(new_n241), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n245), .A2(KEYINPUT30), .A3(new_n240), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n210), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n247), .A2(new_n251), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n254), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT31), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n250), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G472), .A2(G902), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(KEYINPUT32), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT32), .ZN(new_n268));
  INV_X1    g082(.A(new_n250), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n256), .A2(new_n210), .A3(new_n257), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n259), .B1(new_n247), .B2(new_n251), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(new_n254), .A3(KEYINPUT31), .A4(new_n260), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n262), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n266), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n268), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G472), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n248), .A2(new_n249), .A3(new_n198), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n251), .B1(new_n258), .B2(new_n247), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n280), .A2(KEYINPUT29), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n245), .A2(new_n246), .A3(new_n240), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n246), .B1(new_n245), .B2(new_n240), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT28), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n248), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n247), .A2(new_n199), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n251), .A2(KEYINPUT29), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n286), .A2(new_n288), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n282), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n292), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n279), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n278), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT23), .B1(new_n300), .B2(G128), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n238), .A3(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n299), .B1(new_n306), .B2(G110), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n238), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(KEYINPUT24), .A2(G110), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT24), .A2(G110), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT70), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n301), .A2(new_n303), .B1(new_n300), .B2(G128), .ZN(new_n315));
  INV_X1    g129(.A(G110), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n307), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(G146), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n211), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n322), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n211), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n323), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n320), .A2(KEYINPUT72), .A3(G146), .A4(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n306), .A2(G110), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT71), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n315), .A2(KEYINPUT71), .A3(new_n316), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n312), .A2(new_n313), .ZN(new_n336));
  INV_X1    g150(.A(new_n309), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n326), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G137), .ZN(new_n341));
  INV_X1    g155(.A(G953), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(G221), .A3(G234), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n326), .B(new_n344), .C1(new_n332), .C2(new_n339), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n292), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n292), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n350), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n292), .A4(new_n347), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(KEYINPUT74), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n347), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n333), .A2(KEYINPUT71), .B1(new_n336), .B2(new_n337), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n330), .A2(new_n360), .A3(new_n331), .A4(new_n335), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n344), .B1(new_n361), .B2(new_n326), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n353), .A2(G902), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n355), .A2(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n298), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G214), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n234), .A2(new_n239), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n321), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n219), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G224), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G107), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G104), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(KEYINPUT3), .A3(G104), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT3), .B1(new_n377), .B2(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT75), .A3(G101), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(G107), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n378), .B1(new_n388), .B2(new_n380), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n385), .B1(new_n389), .B2(new_n189), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n189), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n384), .A2(new_n390), .A3(KEYINPUT4), .A4(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(G101), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n210), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n207), .A2(KEYINPUT5), .ZN(new_n396));
  INV_X1    g210(.A(G116), .ZN(new_n397));
  OR3_X1    g211(.A1(new_n397), .A2(KEYINPUT5), .A3(G119), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(G113), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n387), .A2(G107), .ZN(new_n402));
  OAI21_X1  g216(.A(G101), .B1(new_n378), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n391), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G122), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n395), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT77), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n395), .B2(new_n405), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(KEYINPUT6), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n412), .B(new_n409), .C1(new_n395), .C2(new_n405), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n376), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n406), .B(KEYINPUT8), .Z(new_n415));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n404), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n373), .A2(new_n418), .A3(new_n375), .ZN(new_n419));
  INV_X1    g233(.A(new_n375), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n371), .A2(new_n372), .B1(KEYINPUT7), .B2(new_n420), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G210), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n425), .A3(new_n423), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n369), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT9), .B(G234), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n292), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n431), .A2(G221), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n292), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n391), .A2(new_n239), .A3(new_n234), .A4(new_n403), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT10), .ZN(new_n436));
  INV_X1    g250(.A(new_n243), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n392), .A2(new_n244), .A3(new_n394), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n342), .A2(G227), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n438), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT10), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n435), .B(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n243), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n404), .A2(new_n370), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n437), .B1(new_n449), .B2(new_n435), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(KEYINPUT12), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(KEYINPUT12), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n439), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n442), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n444), .A2(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n434), .B1(new_n455), .B2(G469), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n451), .A2(new_n452), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n443), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n442), .B1(new_n448), .B2(new_n439), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n433), .B(new_n292), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n432), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n429), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n430), .A2(G217), .A3(new_n342), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT89), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n213), .A2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n238), .A2(G143), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT84), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n221), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(G134), .A3(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n397), .A2(G122), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT81), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT81), .B1(new_n477), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n377), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n397), .A3(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT87), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n478), .B2(G116), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n477), .A2(new_n490), .A3(KEYINPUT14), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .A4(new_n479), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n488), .A2(KEYINPUT85), .B1(G116), .B2(new_n478), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n492), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  OAI21_X1  g310(.A(G107), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT88), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(G107), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n484), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n238), .A2(G143), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n468), .B1(new_n502), .B2(KEYINPUT13), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(KEYINPUT13), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n503), .B2(KEYINPUT82), .ZN(new_n506));
  OAI21_X1  g320(.A(G134), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT83), .B(G134), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  INV_X1    g324(.A(new_n482), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G107), .A3(new_n480), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n512), .A2(new_n483), .B1(new_n221), .B2(new_n473), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n466), .B1(new_n501), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n484), .ZN(new_n516));
  INV_X1    g330(.A(new_n500), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n489), .A2(new_n491), .A3(new_n479), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT86), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n493), .A3(new_n487), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n499), .B1(new_n520), .B2(G107), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n516), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n466), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G478), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT15), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT90), .B(new_n466), .C1(new_n501), .C2(new_n514), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(new_n292), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(KEYINPUT92), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n292), .A3(new_n531), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n527), .A2(KEYINPUT91), .A3(new_n292), .A4(new_n531), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n533), .B1(new_n538), .B2(new_n529), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n540), .B(new_n530), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n319), .B(G146), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT78), .ZN(new_n543));
  INV_X1    g357(.A(G237), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n342), .A3(G214), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n213), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(KEYINPUT18), .A2(G131), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n548), .B(new_n549), .Z(new_n550));
  NOR2_X1   g364(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n548), .B(G131), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT17), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(KEYINPUT17), .A3(G131), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n551), .B1(new_n558), .B2(new_n332), .ZN(new_n559));
  XNOR2_X1  g373(.A(G113), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n387), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n559), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n292), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G475), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT20), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n543), .A2(new_n550), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n319), .B(KEYINPUT19), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n211), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n552), .A2(new_n323), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n571));
  INV_X1    g385(.A(new_n561), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n573), .A3(new_n569), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n559), .A2(new_n561), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n565), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n578), .ZN(new_n580));
  AOI211_X1 g394(.A(KEYINPUT20), .B(new_n580), .C1(new_n575), .C2(new_n576), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n564), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n539), .A2(new_n541), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(G234), .A2(G237), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G952), .A3(new_n342), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT21), .B(G898), .Z(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(G902), .A3(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n464), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n538), .A2(KEYINPUT92), .A3(new_n529), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n561), .B1(new_n570), .B2(KEYINPUT79), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n595), .A2(new_n574), .B1(new_n561), .B2(new_n559), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT20), .B1(new_n596), .B2(new_n580), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n577), .A2(new_n565), .A3(new_n578), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n597), .A2(new_n598), .B1(G475), .B2(new_n563), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n594), .B(new_n599), .C1(new_n600), .C2(new_n533), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(KEYINPUT93), .A3(new_n591), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n367), .B(new_n463), .C1(new_n593), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n527), .A2(new_n605), .A3(new_n531), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n515), .A2(new_n525), .A3(KEYINPUT33), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n528), .A2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n538), .A2(new_n528), .B1(new_n609), .B2(KEYINPUT94), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n606), .A2(new_n607), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n608), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n599), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n429), .A2(new_n592), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n275), .B2(G902), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n275), .B2(new_n276), .ZN(new_n618));
  INV_X1    g432(.A(new_n434), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n453), .A2(new_n454), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n448), .A2(new_n439), .A3(new_n442), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(G469), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n460), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n432), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n366), .A2(new_n618), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n614), .A2(new_n616), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT95), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G6));
  NOR2_X1   g444(.A1(new_n539), .A2(new_n541), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n582), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n616), .A3(new_n626), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT96), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n340), .B(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n355), .A2(new_n358), .B1(new_n364), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n463), .B(new_n640), .C1(new_n593), .C2(new_n602), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT97), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n590), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n586), .B1(new_n646), .B2(KEYINPUT98), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(KEYINPUT98), .B2(new_n646), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT99), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n298), .A2(new_n462), .A3(new_n639), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n632), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  INV_X1    g467(.A(new_n428), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n425), .B1(new_n414), .B2(new_n423), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT38), .Z(new_n657));
  XOR2_X1   g471(.A(new_n649), .B(KEYINPUT39), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n461), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n657), .B1(KEYINPUT40), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(KEYINPUT40), .B2(new_n659), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n582), .B1(new_n539), .B2(new_n541), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n279), .A2(new_n292), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n272), .A2(new_n260), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n242), .A2(new_n247), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n279), .B1(new_n198), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT100), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n278), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n638), .A2(new_n364), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT25), .B1(new_n363), .B2(new_n292), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n674), .B2(new_n354), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n670), .A2(new_n369), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n661), .A2(new_n663), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT101), .B(G143), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G45));
  NAND3_X1  g493(.A1(new_n651), .A2(new_n614), .A3(new_n650), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(new_n292), .B1(new_n458), .B2(new_n459), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n683), .A2(new_n624), .A3(new_n460), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n365), .B(new_n684), .C1(new_n278), .C2(new_n297), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n614), .A3(new_n616), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT102), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT41), .B(G113), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  OAI21_X1  g504(.A(new_n594), .B1(new_n600), .B2(new_n533), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n686), .A2(new_n599), .A3(new_n691), .A4(new_n616), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  AND3_X1   g507(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n292), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT69), .B1(new_n291), .B2(new_n292), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n694), .A2(new_n695), .A3(new_n282), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n277), .B(new_n267), .C1(new_n696), .C2(new_n279), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n368), .B1(new_n654), .B2(new_n655), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n683), .A2(new_n624), .A3(new_n460), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n675), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT93), .B1(new_n601), .B2(new_n591), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n631), .A2(new_n464), .A3(new_n592), .A4(new_n599), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n300), .ZN(G21));
  NAND3_X1  g519(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n198), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n263), .B2(new_n264), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n266), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n365), .A2(new_n617), .A3(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n698), .A2(new_n699), .A3(new_n591), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n691), .A2(new_n710), .A3(new_n582), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  AND3_X1   g527(.A1(new_n675), .A2(new_n617), .A3(new_n709), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n614), .A2(new_n650), .A3(new_n700), .A4(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT103), .B(G125), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G27));
  AOI21_X1  g531(.A(KEYINPUT32), .B1(new_n265), .B2(new_n266), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n275), .A2(new_n268), .A3(new_n276), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n297), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n267), .A2(new_n277), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n427), .A2(new_n368), .A3(new_n428), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n625), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n365), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n538), .A2(new_n528), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n609), .A2(KEYINPUT94), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n613), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n582), .A3(new_n650), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n697), .A2(new_n726), .A3(new_n733), .A4(new_n365), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n228), .ZN(G33));
  OAI211_X1 g551(.A(new_n599), .B(new_n650), .C1(new_n539), .C2(new_n541), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n697), .A2(new_n726), .A3(new_n365), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n221), .ZN(G36));
  NAND2_X1  g555(.A1(new_n730), .A2(new_n599), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT43), .Z(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n618), .A3(new_n675), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n620), .A2(new_n621), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n748), .A2(KEYINPUT105), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT105), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n433), .B1(new_n748), .B2(new_n749), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n746), .B(new_n747), .C1(new_n757), .C2(new_n434), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n434), .B1(new_n754), .B2(new_n755), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT107), .B1(new_n759), .B2(KEYINPUT46), .ZN(new_n760));
  INV_X1    g574(.A(new_n460), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n759), .B2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n624), .A3(new_n658), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n745), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n725), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n744), .B2(KEYINPUT44), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n223), .ZN(G39));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n624), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n763), .A2(new_n772), .A3(new_n624), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n731), .A2(new_n697), .A3(new_n365), .A4(new_n725), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT108), .B(G140), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G42));
  INV_X1    g591(.A(new_n670), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n683), .A2(new_n460), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT49), .Z(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n365), .A3(new_n368), .A4(new_n624), .ZN(new_n781));
  OR4_X1    g595(.A1(new_n778), .A2(new_n781), .A3(new_n657), .A4(new_n742), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n725), .A2(new_n699), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n743), .A2(new_n586), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n297), .B1(new_n278), .B2(KEYINPUT104), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n366), .B1(new_n787), .B2(new_n723), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT48), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(KEYINPUT48), .A3(new_n788), .ZN(new_n792));
  INV_X1    g606(.A(new_n614), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n670), .A2(new_n365), .A3(new_n586), .A4(new_n783), .ZN(new_n794));
  OAI211_X1 g608(.A(G952), .B(new_n342), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n743), .A2(new_n586), .A3(new_n710), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n797), .B2(new_n700), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n610), .A2(new_n599), .A3(new_n613), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n786), .B2(new_n714), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n779), .A2(new_n624), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n771), .B2(new_n773), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n797), .A2(new_n766), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT51), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI22_X1  g621(.A1(new_n803), .A2(new_n807), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n808));
  INV_X1    g622(.A(new_n657), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n369), .A3(new_n684), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n796), .A2(KEYINPUT115), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT115), .B1(new_n796), .B2(new_n810), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(new_n816), .A3(new_n812), .A4(new_n813), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n796), .A2(new_n812), .A3(new_n810), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n799), .B1(new_n808), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n771), .A2(new_n773), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n804), .B1(new_n821), .B2(KEYINPUT114), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(KEYINPUT114), .B2(new_n821), .ZN(new_n823));
  INV_X1    g637(.A(new_n806), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n815), .A2(KEYINPUT117), .A3(new_n817), .A4(new_n818), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(new_n826), .A3(new_n802), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n820), .B1(new_n827), .B2(KEYINPUT51), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n731), .A2(new_n734), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n788), .A2(new_n614), .A3(new_n650), .A4(new_n726), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(KEYINPUT42), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n692), .A2(new_n687), .A3(new_n712), .ZN(new_n833));
  INV_X1    g647(.A(new_n701), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n593), .B2(new_n602), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(KEYINPUT111), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(KEYINPUT53), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n616), .B(new_n626), .C1(new_n632), .C2(new_n614), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n697), .A2(new_n726), .A3(new_n675), .A4(new_n650), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n738), .A2(new_n739), .B1(new_n842), .B2(new_n601), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n730), .A2(new_n582), .A3(new_n650), .A4(new_n714), .ZN(new_n844));
  INV_X1    g658(.A(new_n726), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n603), .A2(new_n641), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT109), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n623), .A2(new_n624), .A3(new_n650), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n675), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n639), .A2(new_n461), .A3(KEYINPUT109), .A4(new_n650), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n670), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n663), .A2(new_n853), .A3(new_n429), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n652), .A2(new_n854), .A3(new_n680), .A4(new_n715), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n650), .B(new_n651), .C1(new_n632), .C2(new_n614), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(KEYINPUT52), .A3(new_n715), .A4(new_n854), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n848), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n829), .B1(new_n840), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n603), .A2(new_n641), .A3(new_n841), .A4(new_n847), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n857), .B2(new_n859), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n692), .A2(new_n687), .A3(new_n712), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n736), .A2(new_n704), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n867), .B2(KEYINPUT111), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n864), .A2(KEYINPUT112), .A3(new_n838), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n848), .A2(new_n860), .A3(new_n867), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n862), .A2(new_n869), .A3(new_n870), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n864), .A2(new_n867), .A3(new_n873), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT113), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n828), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n782), .B1(new_n881), .B2(new_n882), .ZN(G75));
  NAND3_X1  g697(.A1(new_n862), .A2(new_n869), .A3(new_n874), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(G902), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G210), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n411), .A2(new_n413), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(new_n376), .Z(new_n890));
  INV_X1    g704(.A(KEYINPUT55), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(KEYINPUT119), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n888), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n342), .A2(G952), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(KEYINPUT120), .A3(new_n875), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n884), .A2(new_n902), .A3(KEYINPUT54), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n434), .B(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n458), .A2(new_n459), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n903), .A4(new_n904), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n885), .A2(new_n757), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n898), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n913), .A2(new_n596), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n596), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n898), .ZN(G60));
  XNOR2_X1  g730(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n528), .A2(new_n292), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n611), .B1(new_n880), .B2(new_n919), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n611), .A2(new_n901), .A3(new_n903), .A4(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n898), .A3(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT60), .Z(new_n924));
  AOI21_X1  g738(.A(new_n363), .B1(new_n884), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n884), .A2(new_n924), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n898), .B(new_n925), .C1(new_n638), .C2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g742(.A(G953), .B1(new_n588), .B2(new_n374), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n603), .A2(new_n641), .A3(new_n841), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n930), .A2(new_n704), .A3(new_n866), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(G953), .ZN(new_n932));
  INV_X1    g746(.A(G898), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n889), .B1(new_n933), .B2(G953), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n932), .B(new_n934), .Z(G69));
  NAND2_X1  g749(.A1(new_n256), .A2(new_n257), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT123), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n567), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n938), .A2(new_n645), .A3(new_n342), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n663), .A2(new_n788), .A3(new_n429), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n736), .B(new_n740), .C1(new_n764), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n775), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n652), .A2(new_n680), .ZN(new_n944));
  INV_X1    g758(.A(new_n715), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n944), .A2(KEYINPUT124), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT124), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n768), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(KEYINPUT126), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n768), .B2(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n938), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n659), .A2(new_n725), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n367), .B(new_n954), .C1(new_n632), .C2(new_n614), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n765), .B2(new_n767), .ZN(new_n956));
  INV_X1    g770(.A(new_n775), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n946), .A2(new_n677), .A3(new_n947), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n960), .A3(new_n938), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n342), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n940), .B1(new_n953), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n342), .B1(G227), .B2(G900), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n965), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(KEYINPUT125), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(new_n258), .A2(new_n247), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n950), .A2(new_n931), .A3(new_n952), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n664), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n251), .B(new_n970), .C1(new_n971), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n251), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n958), .A2(new_n960), .A3(new_n931), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(new_n974), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n876), .A2(new_n877), .ZN(new_n979));
  INV_X1    g793(.A(new_n281), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n973), .B(new_n979), .C1(new_n980), .C2(new_n665), .ZN(new_n981));
  NOR4_X1   g795(.A1(new_n975), .A2(new_n898), .A3(new_n978), .A4(new_n981), .ZN(G57));
endmodule


