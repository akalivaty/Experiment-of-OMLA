

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U322 ( .A(n319), .B(KEYINPUT17), .ZN(n320) );
  XNOR2_X1 U323 ( .A(n321), .B(n320), .ZN(n323) );
  AND2_X1 U324 ( .A1(G227GAT), .A2(G233GAT), .ZN(n290) );
  NOR2_X1 U325 ( .A1(n477), .A2(n463), .ZN(n464) );
  XNOR2_X1 U326 ( .A(n427), .B(KEYINPUT46), .ZN(n428) );
  XNOR2_X1 U327 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U328 ( .A(n406), .B(n290), .ZN(n324) );
  XNOR2_X1 U329 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n435) );
  XNOR2_X1 U330 ( .A(n364), .B(n324), .ZN(n326) );
  XNOR2_X1 U331 ( .A(n381), .B(n446), .ZN(n382) );
  XNOR2_X1 U332 ( .A(n436), .B(n435), .ZN(n554) );
  XNOR2_X1 U333 ( .A(n346), .B(n332), .ZN(n333) );
  XNOR2_X1 U334 ( .A(n383), .B(n382), .ZN(n426) );
  XNOR2_X1 U335 ( .A(n334), .B(n333), .ZN(n469) );
  XNOR2_X1 U336 ( .A(n488), .B(n487), .ZN(n515) );
  XNOR2_X1 U337 ( .A(n459), .B(G190GAT), .ZN(n460) );
  XNOR2_X1 U338 ( .A(n489), .B(G43GAT), .ZN(n490) );
  XNOR2_X1 U339 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n491), .B(n490), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G92GAT), .B(G99GAT), .Z(n292) );
  XNOR2_X1 U342 ( .A(G29GAT), .B(G106GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n294) );
  XOR2_X1 U344 ( .A(G85GAT), .B(G218GAT), .Z(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n316) );
  INV_X1 U346 ( .A(KEYINPUT79), .ZN(n295) );
  NAND2_X1 U347 ( .A1(G190GAT), .A2(n295), .ZN(n298) );
  INV_X1 U348 ( .A(G190GAT), .ZN(n296) );
  NAND2_X1 U349 ( .A1(n296), .A2(KEYINPUT79), .ZN(n297) );
  NAND2_X1 U350 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U351 ( .A(G162GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U353 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n302) );
  XNOR2_X1 U354 ( .A(KEYINPUT74), .B(KEYINPUT77), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U357 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n306) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(KEYINPUT64), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n310) );
  INV_X1 U361 ( .A(KEYINPUT9), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U363 ( .A(G36GAT), .B(G50GAT), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n414) );
  XNOR2_X1 U366 ( .A(n414), .B(KEYINPUT75), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n318) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n384) );
  INV_X1 U371 ( .A(n384), .ZN(n551) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n321) );
  INV_X1 U373 ( .A(KEYINPUT18), .ZN(n319) );
  XNOR2_X1 U374 ( .A(G190GAT), .B(G183GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n364) );
  XOR2_X1 U376 ( .A(G43GAT), .B(G15GAT), .Z(n406) );
  INV_X1 U377 ( .A(KEYINPUT20), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n334) );
  XNOR2_X1 U379 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n327), .B(KEYINPUT82), .ZN(n328) );
  XOR2_X1 U381 ( .A(n328), .B(KEYINPUT83), .Z(n330) );
  XNOR2_X1 U382 ( .A(G120GAT), .B(G134GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n346) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G71GAT), .ZN(n331) );
  XOR2_X1 U385 ( .A(n331), .B(G176GAT), .Z(n381) );
  XOR2_X1 U386 ( .A(G113GAT), .B(n381), .Z(n332) );
  INV_X1 U387 ( .A(n469), .ZN(n542) );
  XOR2_X1 U388 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n336) );
  XNOR2_X1 U389 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U391 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n350) );
  XNOR2_X1 U393 ( .A(G85GAT), .B(G148GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n339), .B(G57GAT), .ZN(n368) );
  XNOR2_X1 U395 ( .A(G1GAT), .B(G113GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(G29GAT), .B(G141GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n408) );
  INV_X1 U398 ( .A(n408), .ZN(n342) );
  XOR2_X1 U399 ( .A(n368), .B(n342), .Z(n348) );
  XOR2_X1 U400 ( .A(KEYINPUT85), .B(G162GAT), .Z(n344) );
  XNOR2_X1 U401 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(KEYINPUT3), .B(n345), .Z(n456) );
  XNOR2_X1 U404 ( .A(n456), .B(n346), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n352) );
  NAND2_X1 U407 ( .A1(G225GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n476) );
  XNOR2_X1 U409 ( .A(KEYINPUT90), .B(n476), .ZN(n508) );
  INV_X1 U410 ( .A(n508), .ZN(n555) );
  XOR2_X1 U411 ( .A(G92GAT), .B(G64GAT), .Z(n367) );
  XOR2_X1 U412 ( .A(G197GAT), .B(KEYINPUT21), .Z(n354) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n448) );
  XOR2_X1 U415 ( .A(n367), .B(n448), .Z(n356) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U418 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n358) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(KEYINPUT92), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U421 ( .A(n360), .B(n359), .Z(n366) );
  XOR2_X1 U422 ( .A(G176GAT), .B(G204GAT), .Z(n362) );
  XNOR2_X1 U423 ( .A(G36GAT), .B(KEYINPUT78), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n533) );
  XOR2_X1 U427 ( .A(n367), .B(KEYINPUT13), .Z(n370) );
  XNOR2_X1 U428 ( .A(G120GAT), .B(n368), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n372) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U434 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n376) );
  XNOR2_X1 U435 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U437 ( .A(n377), .B(KEYINPUT71), .Z(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U439 ( .A(G106GAT), .B(G78GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n380), .B(G204GAT), .ZN(n446) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT105), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT36), .ZN(n594) );
  XOR2_X1 U443 ( .A(G22GAT), .B(G8GAT), .Z(n418) );
  XOR2_X1 U444 ( .A(G78GAT), .B(G211GAT), .Z(n387) );
  XNOR2_X1 U445 ( .A(G155GAT), .B(G127GAT), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U447 ( .A(n418), .B(n388), .Z(n390) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U450 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n392) );
  XNOR2_X1 U451 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(n394), .B(n393), .Z(n402) );
  XOR2_X1 U454 ( .A(G71GAT), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(G15GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U457 ( .A(KEYINPUT80), .B(G64GAT), .Z(n398) );
  XNOR2_X1 U458 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n577) );
  NOR2_X1 U462 ( .A1(n594), .A2(n577), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n403), .B(KEYINPUT45), .ZN(n423) );
  XOR2_X1 U464 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n405) );
  XNOR2_X1 U465 ( .A(KEYINPUT68), .B(KEYINPUT65), .ZN(n404) );
  XOR2_X1 U466 ( .A(n405), .B(n404), .Z(n422) );
  NAND2_X1 U467 ( .A1(n342), .A2(n406), .ZN(n410) );
  INV_X1 U468 ( .A(n406), .ZN(n407) );
  NAND2_X1 U469 ( .A1(n408), .A2(n407), .ZN(n409) );
  NAND2_X1 U470 ( .A1(n410), .A2(n409), .ZN(n412) );
  AND2_X1 U471 ( .A1(G229GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n413), .B(KEYINPUT66), .ZN(n416) );
  XOR2_X1 U474 ( .A(n414), .B(KEYINPUT29), .Z(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U476 ( .A(G169GAT), .B(n417), .Z(n420) );
  XNOR2_X1 U477 ( .A(n418), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n582) );
  XNOR2_X1 U480 ( .A(n582), .B(KEYINPUT69), .ZN(n569) );
  NAND2_X1 U481 ( .A1(n423), .A2(n569), .ZN(n424) );
  NOR2_X1 U482 ( .A1(n426), .A2(n424), .ZN(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT115), .B(n425), .ZN(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT41), .B(n426), .Z(n560) );
  NAND2_X1 U485 ( .A1(n582), .A2(n560), .ZN(n429) );
  XOR2_X1 U486 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n427) );
  INV_X1 U487 ( .A(n577), .ZN(n588) );
  NOR2_X1 U488 ( .A1(n384), .A2(n588), .ZN(n430) );
  AND2_X1 U489 ( .A1(n431), .A2(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n432), .B(KEYINPUT47), .ZN(n433) );
  AND2_X1 U491 ( .A1(n434), .A2(n433), .ZN(n436) );
  NOR2_X1 U492 ( .A1(n533), .A2(n554), .ZN(n439) );
  XOR2_X1 U493 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n437) );
  XNOR2_X1 U494 ( .A(KEYINPUT122), .B(n437), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U496 ( .A1(n555), .A2(n440), .ZN(n580) );
  XOR2_X1 U497 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n442) );
  XNOR2_X1 U498 ( .A(G141GAT), .B(G22GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U500 ( .A(G50GAT), .B(KEYINPUT74), .Z(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n452) );
  XNOR2_X1 U502 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n445), .B(KEYINPUT23), .ZN(n447) );
  XOR2_X1 U504 ( .A(n447), .B(n446), .Z(n450) );
  XNOR2_X1 U505 ( .A(G148GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n454) );
  NAND2_X1 U508 ( .A1(G228GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n477) );
  NOR2_X1 U511 ( .A1(n580), .A2(n477), .ZN(n457) );
  XOR2_X1 U512 ( .A(KEYINPUT55), .B(n457), .Z(n458) );
  NAND2_X1 U513 ( .A1(n542), .A2(n458), .ZN(n576) );
  NOR2_X1 U514 ( .A1(n551), .A2(n576), .ZN(n461) );
  INV_X1 U515 ( .A(KEYINPUT58), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n426), .A2(n569), .ZN(n496) );
  NOR2_X1 U517 ( .A1(n533), .A2(n469), .ZN(n462) );
  XOR2_X1 U518 ( .A(KEYINPUT97), .B(n462), .Z(n463) );
  NAND2_X1 U519 ( .A1(n464), .A2(KEYINPUT25), .ZN(n468) );
  INV_X1 U520 ( .A(n464), .ZN(n466) );
  INV_X1 U521 ( .A(KEYINPUT25), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n473) );
  XOR2_X1 U524 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n471) );
  NAND2_X1 U525 ( .A1(n469), .A2(n477), .ZN(n470) );
  XOR2_X1 U526 ( .A(n471), .B(n470), .Z(n581) );
  XOR2_X1 U527 ( .A(n533), .B(KEYINPUT94), .Z(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT27), .B(n472), .Z(n478) );
  OR2_X1 U529 ( .A1(n581), .A2(n478), .ZN(n557) );
  NAND2_X1 U530 ( .A1(n473), .A2(n557), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT98), .B(n474), .Z(n475) );
  NOR2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n483) );
  XNOR2_X1 U533 ( .A(KEYINPUT28), .B(n477), .ZN(n514) );
  NOR2_X1 U534 ( .A1(n478), .A2(n514), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n479), .A2(n508), .ZN(n540) );
  XNOR2_X1 U536 ( .A(KEYINPUT84), .B(n542), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n540), .A2(n480), .ZN(n481) );
  XOR2_X1 U538 ( .A(KEYINPUT95), .B(n481), .Z(n482) );
  NOR2_X1 U539 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT99), .B(n484), .Z(n494) );
  NOR2_X1 U541 ( .A1(n594), .A2(n494), .ZN(n485) );
  NAND2_X1 U542 ( .A1(n485), .A2(n577), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n486), .ZN(n530) );
  NAND2_X1 U544 ( .A1(n496), .A2(n530), .ZN(n488) );
  INV_X1 U545 ( .A(KEYINPUT38), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n542), .A2(n515), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n489) );
  NOR2_X1 U548 ( .A1(n384), .A2(n577), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT16), .B(n492), .Z(n493) );
  NOR2_X1 U550 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U551 ( .A(KEYINPUT100), .B(n495), .ZN(n519) );
  NAND2_X1 U552 ( .A1(n496), .A2(n519), .ZN(n505) );
  NOR2_X1 U553 ( .A1(n555), .A2(n505), .ZN(n497) );
  XOR2_X1 U554 ( .A(G1GAT), .B(n497), .Z(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT34), .B(n498), .ZN(G1324GAT) );
  NOR2_X1 U556 ( .A1(n533), .A2(n505), .ZN(n500) );
  XNOR2_X1 U557 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n500), .B(n499), .ZN(G1325GAT) );
  NOR2_X1 U559 ( .A1(n505), .A2(n469), .ZN(n504) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n502) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  INV_X1 U564 ( .A(n514), .ZN(n537) );
  NOR2_X1 U565 ( .A1(n537), .A2(n505), .ZN(n506) );
  XOR2_X1 U566 ( .A(KEYINPUT104), .B(n506), .Z(n507) );
  XNOR2_X1 U567 ( .A(G22GAT), .B(n507), .ZN(G1327GAT) );
  NAND2_X1 U568 ( .A1(n515), .A2(n508), .ZN(n511) );
  XOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .Z(n509) );
  XNOR2_X1 U570 ( .A(KEYINPUT106), .B(n509), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  INV_X1 U572 ( .A(n533), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n512), .A2(n515), .ZN(n513) );
  XNOR2_X1 U574 ( .A(G36GAT), .B(n513), .ZN(G1329GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U576 ( .A(n516), .B(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U577 ( .A(G50GAT), .B(n517), .ZN(G1331GAT) );
  INV_X1 U578 ( .A(n560), .ZN(n573) );
  NOR2_X1 U579 ( .A1(n582), .A2(n573), .ZN(n518) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(n518), .Z(n529) );
  NAND2_X1 U581 ( .A1(n529), .A2(n519), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n555), .A2(n524), .ZN(n520) );
  XOR2_X1 U583 ( .A(n520), .B(KEYINPUT42), .Z(n521) );
  XNOR2_X1 U584 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  NOR2_X1 U585 ( .A1(n533), .A2(n524), .ZN(n522) );
  XOR2_X1 U586 ( .A(G64GAT), .B(n522), .Z(G1333GAT) );
  NOR2_X1 U587 ( .A1(n469), .A2(n524), .ZN(n523) );
  XOR2_X1 U588 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n537), .ZN(n528) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n526) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT111), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U595 ( .A1(n555), .A2(n536), .ZN(n531) );
  XOR2_X1 U596 ( .A(G85GAT), .B(n531), .Z(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT112), .B(n532), .ZN(G1336GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n536), .ZN(n534) );
  XOR2_X1 U599 ( .A(G92GAT), .B(n534), .Z(G1337GAT) );
  NOR2_X1 U600 ( .A1(n469), .A2(n536), .ZN(n535) );
  XOR2_X1 U601 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U605 ( .A1(n554), .A2(n540), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n569), .A2(n550), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  NOR2_X1 U610 ( .A1(n573), .A2(n550), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NOR2_X1 U613 ( .A1(n577), .A2(n550), .ZN(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U616 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XOR2_X1 U620 ( .A(G141GAT), .B(KEYINPUT119), .Z(n559) );
  OR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n582), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1344GAT) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U627 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n588), .A2(n566), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U632 ( .A(G162GAT), .B(KEYINPUT121), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n384), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n576), .ZN(n570) );
  XOR2_X1 U636 ( .A(G169GAT), .B(n570), .Z(G1348GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n573), .A2(n576), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(G1349GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1350GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n584) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n592) );
  NAND2_X1 U647 ( .A1(n592), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U651 ( .A1(n592), .A2(n426), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U654 ( .A1(n592), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(G211GAT), .B(n591), .ZN(G1354GAT) );
  INV_X1 U657 ( .A(n592), .ZN(n593) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(KEYINPUT62), .B(n595), .Z(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

