//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n205), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n205), .B2(new_n207), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT1), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G134gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(G134gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G127gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n217), .B1(new_n221), .B2(new_n215), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n210), .B1(new_n214), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  OR2_X1    g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT24), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  AND2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n228), .B1(new_n227), .B2(new_n231), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(KEYINPUT23), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n235), .A2(KEYINPUT23), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n224), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(G169gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT64), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G169gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT65), .B1(new_n247), .B2(new_n237), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT64), .B(G169gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n242), .ZN(new_n254));
  NOR2_X1   g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n229), .A2(new_n255), .A3(new_n230), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n226), .A2(KEYINPUT24), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n248), .A2(new_n254), .A3(new_n258), .A4(new_n224), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n235), .A2(KEYINPUT26), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(G169gat), .B2(G176gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n236), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n260), .B(new_n226), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n266), .A2(new_n267), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n223), .B1(new_n240), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n227), .A2(new_n231), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n244), .A2(new_n246), .ZN(new_n278));
  INV_X1    g077(.A(new_n242), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n278), .A2(new_n279), .B1(new_n250), .B2(new_n249), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n280), .B2(new_n252), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n251), .B1(new_n253), .B2(new_n242), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT25), .B1(new_n282), .B2(KEYINPUT65), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n269), .B1(new_n266), .B2(new_n267), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n264), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n281), .A2(new_n283), .B1(new_n285), .B2(new_n273), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n203), .A2(new_n208), .A3(new_n209), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n205), .A2(new_n207), .A3(new_n211), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n217), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n209), .B2(KEYINPUT68), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT66), .B1(new_n256), .B2(new_n257), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n239), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT25), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G227gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n202), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G15gat), .B(G43gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(G71gat), .ZN(new_n305));
  INV_X1    g104(.A(G99gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT33), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n240), .A2(new_n275), .A3(new_n223), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n294), .B1(new_n286), .B2(new_n298), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT33), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n301), .B1(new_n276), .B2(new_n299), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n316), .B2(KEYINPUT33), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n315), .A2(new_n317), .A3(new_n307), .A4(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n314), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n303), .B1(new_n322), .B2(KEYINPUT71), .ZN(new_n323));
  INV_X1    g122(.A(new_n307), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT33), .B1(new_n300), .B2(new_n302), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(new_n313), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT72), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n309), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n276), .A2(new_n301), .A3(new_n299), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  INV_X1    g135(.A(new_n309), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n320), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT72), .A3(new_n326), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n336), .B1(new_n340), .B2(KEYINPUT74), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT35), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344));
  INV_X1    g143(.A(G22gat), .ZN(new_n345));
  INV_X1    g144(.A(G228gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G211gat), .B(G218gat), .Z(new_n350));
  AND2_X1   g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(G197gat), .A2(G204gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G211gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G211gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n357), .A3(G218gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n350), .B1(new_n360), .B2(KEYINPUT77), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  INV_X1    g161(.A(new_n350), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT76), .B(G211gat), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT22), .B1(new_n364), .B2(G218gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n362), .B(new_n363), .C1(new_n365), .C2(new_n353), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(G148gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(G148gat), .ZN(new_n374));
  INV_X1    g173(.A(G148gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT82), .A3(G141gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT83), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(KEYINPUT2), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n377), .A2(new_n380), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G141gat), .B(G148gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n383), .B(new_n381), .C1(new_n387), .C2(KEYINPUT2), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n349), .B1(new_n370), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n369), .A3(new_n388), .ZN(new_n391));
  XOR2_X1   g190(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n392));
  AOI22_X1  g191(.A1(new_n391), .A2(new_n392), .B1(new_n361), .B2(new_n366), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT87), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n389), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n368), .B2(new_n369), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398));
  NOR4_X1   g197(.A1(new_n397), .A2(new_n393), .A3(new_n398), .A4(new_n349), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n360), .A2(new_n350), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n392), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n360), .A2(new_n350), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n369), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n389), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n348), .B1(new_n405), .B2(new_n394), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n345), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  NOR4_X1   g207(.A1(new_n395), .A2(new_n399), .A3(new_n406), .A4(G22gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n344), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n394), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  INV_X1    g211(.A(new_n399), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(G22gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n345), .A3(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT88), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n410), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT88), .A4(new_n420), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n342), .A2(new_n343), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  INV_X1    g225(.A(G64gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G92gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n298), .A2(new_n259), .A3(new_n274), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n433), .B2(new_n367), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n433), .B2(new_n432), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n361), .A2(new_n366), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n433), .A2(new_n392), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n431), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n432), .B1(new_n240), .B2(new_n275), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT79), .A3(new_n432), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n445), .A2(new_n448), .A3(new_n441), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n430), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT30), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n450), .A3(new_n430), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n434), .B1(new_n455), .B2(new_n437), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n450), .B1(new_n456), .B2(new_n441), .ZN(new_n457));
  INV_X1    g256(.A(new_n430), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(KEYINPUT81), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n294), .A2(new_n396), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n294), .A2(new_n396), .A3(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n223), .A3(new_n391), .ZN(new_n468));
  NAND2_X1  g267(.A1(G225gat), .A2(G233gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT5), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n465), .A2(new_n466), .A3(new_n468), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(KEYINPUT4), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n223), .B2(new_n389), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n468), .A3(new_n466), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n212), .A2(new_n213), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n222), .B1(new_n477), .B2(new_n289), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n478), .A2(new_n389), .A3(new_n287), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n291), .A2(new_n293), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n480), .A2(new_n210), .B1(new_n388), .B2(new_n386), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n470), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n476), .A2(new_n482), .A3(KEYINPUT5), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n223), .A2(new_n389), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n463), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n488), .B2(new_n470), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(KEYINPUT84), .A3(new_n476), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n473), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G57gat), .B(G85gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n491), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n490), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(new_n501), .B2(new_n472), .ZN(new_n502));
  AOI211_X1 g301(.A(new_n496), .B(new_n473), .C1(new_n485), .C2(new_n490), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n462), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n483), .A2(new_n484), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT84), .B1(new_n489), .B2(new_n476), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n472), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n496), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n497), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n499), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n505), .B2(new_n513), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n328), .A2(new_n336), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n340), .A2(new_n334), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n453), .A2(new_n454), .A3(new_n461), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n422), .A2(new_n423), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n515), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n425), .A2(new_n506), .B1(new_n521), .B2(new_n343), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n470), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n524), .B(KEYINPUT39), .C1(new_n470), .C2(new_n488), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n497), .C1(KEYINPUT39), .C2(new_n524), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT89), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n526), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n462), .A2(new_n529), .A3(new_n510), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n443), .A2(KEYINPUT37), .A3(new_n450), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n457), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n533), .A3(new_n430), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n451), .B1(new_n534), .B2(KEYINPUT38), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n535), .B(new_n514), .C1(new_n505), .C2(new_n513), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT38), .B(new_n458), .C1(new_n457), .C2(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n440), .A2(KEYINPUT91), .A3(new_n441), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(new_n456), .B2(new_n442), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n445), .A2(new_n448), .A3(new_n442), .A4(new_n449), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT37), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT92), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n537), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n520), .B(new_n530), .C1(new_n536), .C2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n335), .A2(new_n341), .A3(KEYINPUT36), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT75), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n516), .A2(new_n552), .A3(new_n517), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n506), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n424), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n335), .A2(new_n341), .A3(KEYINPUT75), .A4(KEYINPUT36), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(new_n554), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n522), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  OR2_X1    g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G57gat), .B(G64gat), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT97), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n560), .A3(new_n561), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(G1gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G1gat), .B2(new_n571), .ZN(new_n574));
  INV_X1    g373(.A(G8gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT98), .ZN(new_n578));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G183gat), .B(G211gat), .Z(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  INV_X1    g389(.A(G106gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT8), .B1(new_n306), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n590), .B(new_n592), .C1(G85gat), .C2(G92gat), .ZN(new_n593));
  XOR2_X1   g392(.A(G99gat), .B(G106gat), .Z(new_n594));
  OR3_X1    g393(.A1(new_n593), .A2(KEYINPUT99), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT99), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT100), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n599), .A3(new_n596), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n598), .A2(new_n600), .B1(new_n594), .B2(new_n593), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G29gat), .ZN(new_n603));
  INV_X1    g402(.A(G36gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT14), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT14), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(G29gat), .B2(G36gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G43gat), .B(G50gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT15), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT15), .ZN(new_n614));
  NAND2_X1  g413(.A1(G29gat), .A2(G36gat), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n610), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n608), .A2(KEYINPUT93), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n608), .B2(KEYINPUT93), .ZN(new_n618));
  OAI211_X1 g417(.A(KEYINPUT15), .B(new_n611), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT17), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n602), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n620), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n602), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n622), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n622), .B2(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n628), .B2(KEYINPUT101), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n631), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n588), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n559), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n576), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n624), .A2(new_n576), .ZN(new_n642));
  NAND2_X1  g441(.A1(G229gat), .A2(G233gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT18), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n620), .B(new_n576), .Z(new_n647));
  XOR2_X1   g446(.A(new_n643), .B(KEYINPUT13), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT11), .B(G169gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G197gat), .ZN(new_n653));
  XOR2_X1   g452(.A(G113gat), .B(G141gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n646), .A2(new_n656), .A3(new_n649), .A4(new_n650), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n593), .A2(new_n594), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n569), .A2(new_n597), .A3(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n665), .B(new_n667), .C1(new_n601), .C2(new_n569), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n601), .A2(KEYINPUT102), .A3(KEYINPUT10), .A4(new_n569), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G176gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G204gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n667), .B1(new_n601), .B2(new_n569), .ZN(new_n676));
  INV_X1    g475(.A(new_n671), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n672), .B(new_n680), .C1(new_n679), .C2(new_n678), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n672), .A2(new_n678), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n675), .B(KEYINPUT104), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n661), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n638), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n505), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n687), .B(new_n462), .C1(KEYINPUT16), .C2(G8gat), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n572), .A2(new_n575), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n575), .B1(new_n687), .B2(new_n462), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(G1325gat));
  AND2_X1   g498(.A1(new_n554), .A2(new_n557), .ZN(new_n700));
  OAI21_X1  g499(.A(G15gat), .B1(new_n686), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n687), .A2(new_n518), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(G15gat), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT106), .Z(G1326gat));
  NOR2_X1   g503(.A1(new_n686), .A2(new_n520), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(new_n636), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n522), .B2(new_n558), .ZN(new_n709));
  INV_X1    g508(.A(new_n588), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n661), .A3(new_n684), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n603), .A3(new_n505), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n335), .A2(new_n341), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(KEYINPUT35), .A3(new_n506), .A4(new_n520), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n340), .A2(new_n334), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n337), .B(new_n336), .C1(new_n338), .C2(new_n339), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n423), .B(new_n422), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n500), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n513), .B1(new_n512), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT90), .B1(new_n504), .B2(new_n499), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n519), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n343), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n717), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n722), .A2(new_n723), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(new_n535), .A3(new_n545), .A4(new_n547), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n530), .A2(new_n520), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n728), .A2(new_n729), .B1(new_n555), .B2(new_n424), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n700), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n731), .B2(new_n708), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n709), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n711), .B(KEYINPUT107), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n505), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n715), .A2(new_n739), .ZN(G1328gat));
  NAND3_X1  g539(.A1(new_n713), .A2(new_n604), .A3(new_n462), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT108), .ZN(new_n745));
  OAI21_X1  g544(.A(G36gat), .B1(new_n737), .B2(new_n519), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n745), .B(new_n746), .C1(new_n743), .C2(new_n742), .ZN(G1329gat));
  OAI21_X1  g546(.A(G43gat), .B1(new_n737), .B2(new_n700), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT47), .B1(new_n748), .B2(KEYINPUT109), .ZN(new_n749));
  INV_X1    g548(.A(G43gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n713), .A2(new_n750), .A3(new_n518), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n749), .B(new_n752), .ZN(G1330gat));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n424), .A3(new_n736), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(G50gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n712), .A2(G50gat), .A3(new_n520), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g557(.A1(new_n638), .A2(new_n661), .A3(new_n684), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n505), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT111), .B(G57gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1332gat));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n759), .B(new_n462), .C1(new_n763), .C2(new_n427), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n427), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(new_n700), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G71gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n759), .A2(new_n518), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(G71gat), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g571(.A1(new_n759), .A2(new_n424), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n661), .A2(new_n588), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT112), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n559), .B2(new_n636), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT114), .B(new_n708), .C1(new_n522), .C2(new_n558), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT51), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n783), .A2(KEYINPUT115), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n505), .A4(new_n684), .ZN(new_n786));
  INV_X1    g585(.A(G85gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n709), .A2(new_n733), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT44), .B(new_n708), .C1(new_n522), .C2(new_n558), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n684), .B(new_n776), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n735), .A2(KEYINPUT113), .A3(new_n684), .A4(new_n776), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n786), .A2(new_n787), .B1(new_n505), .B2(new_n794), .ZN(G1336gat));
  NAND3_X1  g594(.A1(new_n684), .A2(new_n429), .A3(new_n462), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT116), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n784), .A2(new_n785), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  OAI21_X1  g599(.A(G92gat), .B1(new_n790), .B2(new_n519), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n792), .A2(new_n793), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n429), .B1(new_n803), .B2(new_n462), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n782), .A2(new_n783), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n798), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT117), .B(new_n797), .C1(new_n782), .C2(new_n783), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n804), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n802), .B1(new_n809), .B2(new_n800), .ZN(G1337gat));
  AOI211_X1 g609(.A(new_n306), .B(new_n700), .C1(new_n792), .C2(new_n793), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n784), .A2(new_n785), .A3(new_n684), .A4(new_n518), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n306), .B2(new_n812), .ZN(G1338gat));
  AOI21_X1  g612(.A(new_n591), .B1(new_n803), .B2(new_n424), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n520), .A2(G106gat), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n806), .A2(new_n684), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT53), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n784), .A2(new_n785), .A3(new_n684), .A4(new_n815), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  OAI21_X1  g618(.A(G106gat), .B1(new_n790), .B2(new_n520), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(G1339gat));
  NAND4_X1  g621(.A1(new_n664), .A2(new_n668), .A3(new_n677), .A4(new_n669), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n672), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g623(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n825));
  NAND3_X1  g624(.A1(new_n670), .A2(new_n671), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n675), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n681), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n660), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n643), .B1(new_n641), .B2(new_n642), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n647), .A2(new_n648), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n655), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n659), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n636), .B1(new_n837), .B2(new_n684), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n831), .A2(new_n837), .A3(new_n832), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n636), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n841), .A3(new_n588), .ZN(new_n842));
  INV_X1    g641(.A(new_n684), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n637), .A2(new_n661), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n738), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n342), .A2(new_n424), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n519), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n206), .A3(new_n660), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n720), .B1(new_n842), .B2(new_n844), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n738), .A2(new_n462), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n661), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT119), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n852), .B2(new_n843), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n843), .A2(new_n462), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n845), .A2(new_n204), .A3(new_n846), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1341gat));
  NOR3_X1   g658(.A1(new_n852), .A2(new_n216), .A3(new_n588), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n848), .A2(new_n710), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n216), .ZN(G1342gat));
  NOR3_X1   g661(.A1(new_n847), .A2(G134gat), .A3(new_n708), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n852), .B2(new_n708), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT120), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(G1343gat));
  AOI21_X1  g668(.A(new_n520), .B1(new_n842), .B2(new_n844), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n700), .A2(new_n851), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G141gat), .A3(new_n661), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n876), .B(new_n520), .C1(new_n842), .C2(new_n844), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n660), .B(new_n872), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n878), .B2(G141gat), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT58), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  AOI221_X4 g682(.A(new_n874), .B1(new_n880), .B2(new_n883), .C1(G141gat), .C2(new_n878), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n767), .A2(new_n520), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n845), .A2(new_n375), .A3(new_n857), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n842), .A2(new_n844), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n876), .B1(new_n888), .B2(new_n520), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n684), .A3(new_n872), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(G148gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n892), .B2(G148gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(G1345gat));
  INV_X1    g695(.A(G155gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n873), .B2(new_n588), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n891), .A2(new_n872), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n588), .A2(new_n897), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT122), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(G1346gat));
  INV_X1    g703(.A(new_n873), .ZN(new_n905));
  AOI21_X1  g704(.A(G162gat), .B1(new_n905), .B2(new_n636), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n899), .A2(new_n708), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n519), .A2(new_n505), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n850), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n661), .ZN(new_n911));
  AOI211_X1 g710(.A(new_n505), .B(new_n519), .C1(new_n842), .C2(new_n844), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n846), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n660), .A2(new_n278), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1348gat));
  NOR3_X1   g714(.A1(new_n910), .A2(new_n241), .A3(new_n843), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n684), .A3(new_n846), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n241), .B2(new_n917), .ZN(G1349gat));
  OAI21_X1  g717(.A(G183gat), .B1(new_n910), .B2(new_n588), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n710), .A2(new_n266), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g721(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n923));
  OAI211_X1 g722(.A(G190gat), .B(new_n923), .C1(new_n910), .C2(new_n708), .ZN(new_n924));
  NOR2_X1   g723(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n912), .A2(new_n267), .A3(new_n846), .A4(new_n636), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G1351gat));
  NAND2_X1  g728(.A1(new_n700), .A2(new_n909), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT125), .Z(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n889), .B2(new_n890), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n661), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n886), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(G197gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n661), .B2(new_n936), .ZN(G1352gat));
  XOR2_X1   g736(.A(KEYINPUT126), .B(G204gat), .Z(new_n938));
  OR3_X1    g737(.A1(new_n935), .A2(new_n843), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n891), .A2(new_n684), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n938), .B1(new_n944), .B2(new_n931), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n943), .B(new_n945), .C1(new_n941), .C2(new_n939), .ZN(G1353gat));
  OR3_X1    g745(.A1(new_n935), .A2(new_n364), .A3(new_n588), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n710), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  OAI21_X1  g750(.A(G218gat), .B1(new_n933), .B2(new_n708), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n935), .A2(G218gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n708), .B2(new_n953), .ZN(G1355gat));
endmodule


