//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G226), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n202), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR4_X1   g0020(.A1(new_n209), .A2(new_n214), .A3(new_n217), .A4(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT65), .B(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G116), .ZN(new_n224));
  INV_X1    g0024(.A(G270), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G1), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n219), .B(new_n234), .C1(new_n211), .C2(new_n213), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n236), .A2(new_n228), .ZN(new_n237));
  OAI21_X1  g0037(.A(G50), .B1(G58), .B2(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT64), .ZN(new_n239));
  AOI22_X1  g0039(.A1(new_n235), .A2(KEYINPUT0), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  OAI211_X1 g0040(.A(new_n232), .B(new_n240), .C1(KEYINPUT0), .C2(new_n235), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n216), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT2), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n206), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G264), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n225), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(G107), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(new_n224), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  INV_X1    g0057(.A(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT10), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n258), .A2(KEYINPUT10), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n227), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G222), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(new_n269), .B1(G223), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n272), .B1(new_n269), .B2(new_n268), .C1(new_n207), .C2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n236), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n263), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n276), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(new_n261), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(G190), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n277), .A2(new_n280), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT71), .B(G200), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n228), .A2(G1), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT68), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n202), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(new_n228), .A3(G1), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n236), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(KEYINPUT67), .A3(new_n236), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n203), .A2(G20), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G150), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n298), .B(new_n300), .C1(new_n301), .C2(new_n304), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n291), .A2(KEYINPUT67), .A3(new_n236), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT67), .B1(new_n291), .B2(new_n236), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n305), .A2(new_n308), .B1(new_n202), .B2(new_n290), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT9), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n259), .B(new_n260), .C1(new_n285), .C2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n284), .B1(new_n277), .B2(new_n280), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G190), .B2(new_n282), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n315), .A2(new_n258), .A3(KEYINPUT10), .A4(new_n311), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n282), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n310), .C1(G169), .C2(new_n282), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n279), .A2(G238), .ZN(new_n321));
  INV_X1    g0121(.A(new_n263), .ZN(new_n322));
  AND3_X1   g0122(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n266), .B1(new_n216), .B2(G1698), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n206), .A2(new_n270), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n321), .B(new_n322), .C1(new_n328), .C2(new_n278), .ZN(new_n329));
  XOR2_X1   g0129(.A(new_n329), .B(KEYINPUT13), .Z(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT14), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(G179), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n329), .B(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(G169), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n287), .A2(new_n290), .A3(new_n292), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G68), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n303), .A2(G77), .B1(new_n299), .B2(G50), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n228), .B2(G68), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT11), .A3(new_n308), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n286), .A2(G13), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(G68), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT11), .B1(new_n341), .B2(new_n308), .ZN(new_n347));
  OR3_X1    g0147(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n334), .B2(G200), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n330), .A2(G190), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n299), .B(KEYINPUT69), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n353), .A2(new_n301), .B1(new_n228), .B2(new_n207), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT70), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT15), .B(G87), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n304), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n292), .B1(new_n207), .B2(new_n290), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n338), .A2(G77), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n267), .A2(G232), .ZN(new_n362));
  INV_X1    g0162(.A(new_n271), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n362), .B1(new_n212), .B2(new_n273), .C1(new_n363), .C2(new_n223), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n263), .B1(new_n364), .B2(new_n276), .ZN(new_n365));
  INV_X1    g0165(.A(new_n279), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n208), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n331), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n367), .A2(G179), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n349), .A2(new_n352), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n320), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(G223), .B(new_n270), .C1(new_n264), .C2(new_n265), .ZN(new_n373));
  OAI211_X1 g0173(.A(G226), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT76), .A4(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n276), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n263), .B1(new_n279), .B2(G232), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n382), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT78), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n380), .A2(new_n388), .A3(new_n381), .A4(new_n382), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n287), .A2(new_n301), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n296), .B1(new_n290), .B2(new_n301), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n273), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n266), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n228), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(G68), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n215), .A2(new_n222), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n201), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n299), .A2(KEYINPUT74), .A3(G159), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT74), .B1(new_n299), .B2(G159), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n394), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n292), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n222), .B1(new_n396), .B2(new_n397), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n406), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n393), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n390), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT79), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT79), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n416), .A3(KEYINPUT17), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n390), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT80), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT80), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n390), .A2(new_n412), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n415), .A2(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n412), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n380), .A2(new_n317), .A3(new_n382), .ZN(new_n425));
  AOI21_X1  g0225(.A(G169), .B1(new_n380), .B2(new_n382), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT77), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n385), .B2(G179), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT18), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n367), .A2(new_n381), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n367), .A2(new_n283), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n433), .A2(new_n359), .A3(new_n360), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n372), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(G244), .B(new_n270), .C1(new_n264), .C2(new_n265), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n438), .A2(new_n208), .A3(G1698), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n219), .A2(new_n270), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n273), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n276), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(G274), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n276), .B1(new_n448), .B2(new_n446), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G257), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n386), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n445), .A2(new_n452), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n453), .A2(new_n454), .B1(new_n455), .B2(new_n381), .ZN(new_n456));
  INV_X1    g0256(.A(new_n455), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT82), .A3(G190), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT81), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n227), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n296), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n344), .B(new_n461), .C1(new_n306), .C2(new_n307), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n210), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n399), .A2(G107), .A3(new_n400), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n299), .A2(G77), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n212), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n210), .A2(new_n212), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G20), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n466), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n465), .B1(new_n474), .B2(new_n292), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n344), .A2(G97), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT83), .B1(new_n459), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n455), .A2(G179), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n478), .B(new_n481), .C1(G169), .C2(new_n457), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n476), .B(new_n465), .C1(new_n474), .C2(new_n292), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n458), .A4(new_n456), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n227), .A2(G45), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(G250), .C1(new_n275), .C2(new_n236), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n448), .A2(G274), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT84), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n495));
  OAI211_X1 g0295(.A(G238), .B(new_n270), .C1(new_n264), .C2(new_n265), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n302), .C2(new_n224), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n276), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n494), .A2(KEYINPUT85), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT85), .B1(new_n494), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(G190), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT19), .B1(new_n323), .B2(new_n324), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n228), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n273), .A2(new_n228), .A3(G68), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT19), .B1(new_n303), .B2(G97), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n510), .A2(new_n408), .B1(new_n344), .B2(new_n356), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n460), .B1(new_n296), .B2(new_n461), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n513));
  OAI21_X1  g0313(.A(G87), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT86), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n462), .A2(new_n464), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(G87), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n511), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n500), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n494), .A2(KEYINPUT85), .A3(new_n498), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n283), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT87), .B(G190), .C1(new_n499), .C2(new_n500), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n503), .A2(new_n519), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n521), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n317), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n331), .A3(new_n521), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n357), .B1(new_n462), .B2(new_n464), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n511), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT92), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n273), .A2(G250), .A3(new_n270), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G294), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n450), .B1(new_n536), .B2(new_n276), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n451), .A2(G264), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n537), .A2(G179), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n331), .B1(new_n537), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n532), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G169), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(G179), .A3(new_n538), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(KEYINPUT92), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT91), .B1(new_n212), .B2(G20), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(G116), .B2(new_n303), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n228), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT89), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT90), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT90), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(new_n558), .A3(new_n554), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n551), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT24), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n552), .A2(new_n558), .A3(new_n554), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(new_n552), .B2(new_n554), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n553), .B(KEYINPUT22), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n551), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n408), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n212), .B1(new_n462), .B2(new_n464), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n290), .A2(new_n212), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT25), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n546), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n408), .A2(new_n344), .A3(G116), .A4(new_n461), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n443), .B(new_n228), .C1(G33), .C2(new_n210), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n292), .C1(new_n228), .C2(G116), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT20), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  OAI221_X1 g0383(.A(new_n578), .B1(G116), .B2(new_n344), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n225), .B(new_n276), .C1(new_n448), .C2(new_n446), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n266), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n270), .A2(G257), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G264), .A2(G1698), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n264), .C2(new_n265), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n276), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT88), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n587), .A2(KEYINPUT88), .A3(new_n276), .A4(new_n590), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n585), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n584), .A2(G179), .A3(new_n449), .A4(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n331), .B1(new_n595), .B2(new_n449), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n584), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n601), .A3(new_n584), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n597), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n569), .B1(new_n568), .B2(new_n551), .ZN(new_n604));
  INV_X1    g0404(.A(new_n551), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT24), .B(new_n605), .C1(new_n566), .C2(new_n567), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n292), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n542), .A2(new_n386), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G190), .B2(new_n542), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n609), .A3(new_n575), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n595), .A2(new_n449), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G200), .ZN(new_n612));
  INV_X1    g0412(.A(new_n584), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n381), .C2(new_n611), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n577), .A2(new_n603), .A3(new_n610), .A4(new_n614), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n436), .A2(new_n486), .A3(new_n531), .A4(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n436), .ZN(new_n617));
  AOI21_X1  g0417(.A(G169), .B1(new_n445), .B2(new_n452), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n618), .B(new_n480), .C1(new_n475), .C2(new_n477), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n524), .A2(new_n619), .A3(new_n530), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n494), .A2(new_n498), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n331), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n526), .A2(new_n529), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n283), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n503), .A2(new_n519), .A3(new_n523), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n539), .A2(new_n540), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n607), .B2(new_n575), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n601), .A2(new_n611), .A3(G169), .A4(new_n584), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n601), .B1(new_n598), .B2(new_n584), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n596), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n624), .B(new_n626), .C1(new_n628), .C2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n610), .A2(new_n479), .A3(new_n482), .A4(new_n485), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n621), .B(new_n624), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n624), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n635), .A2(KEYINPUT26), .A3(new_n482), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n617), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n319), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT18), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n430), .B(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n370), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n352), .B1(new_n337), .B2(new_n348), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n423), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n313), .A2(new_n316), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT93), .Z(G369));
  NOR2_X1   g0448(.A1(new_n289), .A2(G20), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n227), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n613), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n614), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n631), .A2(new_n659), .A3(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(KEYINPUT94), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(KEYINPUT94), .B2(new_n658), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n577), .A2(new_n656), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n577), .A2(new_n610), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n655), .B1(new_n571), .B2(new_n576), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n631), .A3(new_n656), .ZN(new_n670));
  INV_X1    g0470(.A(new_n628), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n655), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n669), .A2(new_n672), .ZN(G399));
  NOR2_X1   g0473(.A1(new_n234), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n504), .A2(new_n224), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(G1), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n239), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n675), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n637), .A2(new_n656), .ZN(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n685));
  INV_X1    g0485(.A(new_n635), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n577), .A2(new_n603), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n685), .B(new_n624), .C1(new_n688), .C2(new_n633), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n686), .B2(new_n619), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT29), .B(new_n656), .C1(new_n689), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n595), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n544), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT95), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n455), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n525), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n696), .B2(new_n697), .ZN(new_n700));
  AOI21_X1  g0500(.A(G179), .B1(new_n537), .B2(new_n538), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n611), .A2(new_n701), .A3(new_n455), .A4(new_n622), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n696), .A2(new_n697), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n525), .A2(new_n695), .A3(new_n703), .A4(new_n698), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n655), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AND4_X1   g0507(.A1(new_n577), .A2(new_n603), .A3(new_n610), .A4(new_n614), .ZN(new_n708));
  INV_X1    g0508(.A(new_n486), .ZN(new_n709));
  INV_X1    g0509(.A(new_n531), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n656), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n707), .B1(new_n711), .B2(KEYINPUT31), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(G330), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n693), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n681), .B1(new_n716), .B2(G1), .ZN(G364));
  NAND2_X1  g0517(.A1(new_n649), .A2(G45), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n675), .A2(G1), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n663), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n662), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n253), .A2(G45), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n234), .A2(new_n273), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n723), .B(new_n724), .C1(G45), .C2(new_n679), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n233), .A2(G355), .A3(new_n273), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n725), .B(new_n726), .C1(G116), .C2(new_n233), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n236), .B1(G20), .B2(new_n331), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n719), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT97), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n228), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n283), .A2(G190), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n218), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n283), .A2(new_n381), .A3(new_n735), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n212), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n381), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n317), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G97), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n228), .A2(new_n317), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n381), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G50), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n740), .A2(new_n273), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT98), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT98), .B1(new_n228), .B2(new_n317), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n751), .A2(new_n741), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n754), .A2(new_n215), .B1(new_n207), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n745), .A2(new_n381), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n222), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n735), .A2(new_n755), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n749), .A2(new_n757), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n754), .A2(new_n766), .B1(new_n767), .B2(new_n756), .ZN(new_n768));
  INV_X1    g0568(.A(new_n758), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n273), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n747), .A2(G326), .ZN(new_n772));
  INV_X1    g0572(.A(new_n760), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G329), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n743), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n779), .A2(new_n738), .B1(new_n736), .B2(new_n586), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n768), .A2(new_n775), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n731), .B1(new_n765), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n730), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n734), .B(new_n782), .C1(new_n662), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n722), .A2(new_n784), .ZN(G396));
  AND4_X1   g0585(.A1(new_n361), .A2(new_n368), .A3(new_n369), .A4(new_n656), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n361), .A2(new_n655), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n435), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n788), .B2(new_n370), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n682), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n656), .B(new_n789), .C1(new_n634), .C2(new_n636), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(new_n715), .Z(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n719), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n731), .A2(new_n728), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n207), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G303), .A2(new_n747), .B1(new_n769), .B2(G283), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n273), .B1(new_n773), .B2(G311), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n798), .A2(new_n744), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n736), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G107), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n738), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G87), .ZN(new_n804));
  INV_X1    g0604(.A(new_n756), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G116), .A2(new_n805), .B1(new_n753), .B2(G294), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT100), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n738), .A2(new_n222), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n273), .B1(new_n736), .B2(new_n202), .C1(new_n776), .C2(new_n215), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n805), .A2(G159), .B1(G137), .B2(new_n747), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n753), .A2(G143), .ZN(new_n812));
  INV_X1    g0612(.A(G150), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n758), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT34), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n809), .B(new_n810), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n815), .B2(new_n814), .C1(new_n817), .C2(new_n760), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n808), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n719), .B1(new_n819), .B2(new_n731), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n797), .B(new_n820), .C1(new_n789), .C2(new_n729), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n795), .A2(new_n821), .ZN(G384));
  NAND2_X1  g0622(.A1(new_n431), .A2(new_n653), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n394), .B1(new_n409), .B2(new_n406), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n824), .A2(new_n308), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n392), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n427), .A2(new_n827), .A3(new_n429), .ZN(new_n828));
  INV_X1    g0628(.A(new_n653), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n828), .A2(new_n413), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n424), .A2(new_n829), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n430), .A2(new_n833), .A3(new_n413), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n832), .A2(KEYINPUT103), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT103), .B1(new_n832), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n420), .A2(new_n422), .ZN(new_n839));
  AOI211_X1 g0639(.A(KEYINPUT79), .B(new_n418), .C1(new_n390), .C2(new_n412), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n416), .B1(new_n413), .B2(KEYINPUT17), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n830), .B1(new_n842), .B2(new_n641), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n838), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n832), .A2(new_n835), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n832), .A2(new_n835), .A3(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n830), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n423), .B2(new_n431), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n786), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n792), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n348), .A2(new_n655), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n349), .A2(new_n352), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n352), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n348), .B(new_n655), .C1(new_n859), .C2(new_n337), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n854), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n850), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n833), .B1(new_n842), .B2(new_n641), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n430), .A2(new_n413), .A3(new_n833), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(new_n834), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n844), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT39), .B1(new_n845), .B2(new_n853), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n844), .B1(new_n838), .B2(new_n843), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n865), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n349), .A2(new_n655), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n823), .B(new_n864), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n684), .A2(new_n617), .A3(new_n692), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n646), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n882), .B(new_n884), .Z(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n713), .B(KEYINPUT106), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n789), .B(new_n861), .C1(new_n712), .C2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n854), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n712), .A2(new_n887), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n858), .A2(new_n860), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n790), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n870), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n436), .A2(new_n890), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n885), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n227), .B2(new_n649), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n224), .B1(new_n472), .B2(KEYINPUT35), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n237), .C1(KEYINPUT35), .C2(new_n472), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT36), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n679), .A2(new_n207), .A3(new_n402), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n202), .B2(G68), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n905), .A2(new_n227), .A3(G13), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT101), .Z(new_n907));
  NAND3_X1  g0707(.A1(new_n900), .A2(new_n903), .A3(new_n907), .ZN(G367));
  OR2_X1    g0708(.A1(new_n519), .A2(new_n656), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n686), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n624), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n709), .B1(new_n483), .B2(new_n656), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n670), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  OR2_X1    g0715(.A1(new_n913), .A2(new_n577), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n655), .B1(new_n916), .B2(new_n482), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n912), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n619), .A2(new_n655), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n664), .A2(new_n668), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n918), .B(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n674), .B(KEYINPUT41), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n668), .B1(new_n603), .B2(new_n655), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT108), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n670), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(new_n663), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT109), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n930), .A2(new_n931), .A3(new_n716), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n930), .B2(new_n716), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n920), .A2(new_n672), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT44), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n920), .A2(new_n672), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n669), .A2(KEYINPUT107), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n926), .B1(new_n942), .B2(new_n716), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n718), .A2(G1), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n924), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n736), .B2(new_n224), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(new_n754), .C2(new_n586), .ZN(new_n949));
  INV_X1    g0749(.A(new_n747), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n950), .A2(new_n767), .B1(new_n776), .B2(new_n212), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n273), .B(new_n951), .C1(G294), .C2(new_n769), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n773), .A2(G317), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n210), .C2(new_n738), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n949), .B(new_n954), .C1(G283), .C2(new_n805), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n753), .A2(G150), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n803), .A2(G77), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n743), .A2(G68), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(new_n215), .C2(new_n736), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G143), .A2(new_n747), .B1(new_n769), .B2(G159), .ZN(new_n960));
  INV_X1    g0760(.A(G137), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n273), .C1(new_n961), .C2(new_n760), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n959), .B(new_n962), .C1(G50), .C2(new_n805), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n955), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  AOI21_X1  g0765(.A(new_n719), .B1(new_n965), .B2(new_n731), .ZN(new_n966));
  INV_X1    g0766(.A(new_n724), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n732), .B1(new_n233), .B2(new_n357), .C1(new_n249), .C2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT110), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n966), .B(new_n969), .C1(new_n911), .C2(new_n783), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n945), .A2(new_n970), .ZN(G387));
  AOI22_X1  g0771(.A1(G303), .A2(new_n805), .B1(new_n753), .B2(G317), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n972), .A2(KEYINPUT111), .B1(G311), .B2(new_n769), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(KEYINPUT111), .B2(new_n972), .C1(new_n766), .C2(new_n950), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n779), .B2(new_n776), .C1(new_n777), .C2(new_n736), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT49), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n773), .A2(G326), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n273), .B1(new_n803), .B2(G116), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n776), .A2(new_n357), .B1(new_n301), .B2(new_n758), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n266), .B(new_n983), .C1(G159), .C2(new_n747), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n773), .A2(G150), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G68), .A2(new_n805), .B1(new_n753), .B2(G50), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G77), .A2(new_n801), .B1(new_n803), .B2(G97), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n731), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n301), .A2(G50), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT50), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n677), .B1(new_n222), .B2(new_n207), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AOI211_X1 g0793(.A(G45), .B(new_n993), .C1(new_n992), .C2(new_n991), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n724), .B1(new_n246), .B2(new_n447), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n233), .A2(new_n273), .A3(new_n676), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n233), .A2(G107), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n732), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n990), .A2(new_n720), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT112), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n668), .B2(new_n730), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n944), .B2(new_n930), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n674), .B1(new_n716), .B2(new_n930), .C1(new_n932), .C2(new_n933), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(G393));
  OAI21_X1  g0805(.A(new_n939), .B1(KEYINPUT113), .B2(new_n669), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n669), .A2(KEYINPUT113), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  OAI211_X1 g0808(.A(new_n942), .B(new_n674), .C1(new_n934), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n920), .A2(new_n730), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n776), .A2(new_n207), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G50), .B2(new_n769), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n266), .B1(new_n773), .B2(G143), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n804), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n301), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n805), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n753), .A2(G159), .B1(G150), .B2(new_n747), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT51), .Z(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(new_n222), .C2(new_n736), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT114), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n266), .B1(new_n756), .B2(new_n777), .C1(new_n776), .C2(new_n224), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n739), .B(new_n1021), .C1(G303), .C2(new_n769), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n753), .A2(G311), .B1(G317), .B2(new_n747), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT52), .Z(new_n1024));
  OAI22_X1  g0824(.A1(new_n736), .A2(new_n779), .B1(new_n766), .B2(new_n760), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT115), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n719), .B1(new_n1028), .B2(new_n731), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n732), .B1(new_n210), .B2(new_n233), .C1(new_n256), .C2(new_n967), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1010), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1008), .B2(new_n944), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1009), .A2(new_n1032), .ZN(G390));
  NAND2_X1  g0833(.A1(new_n789), .A2(G330), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n615), .A2(new_n486), .A3(new_n531), .A4(new_n655), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT31), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n706), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1034), .B1(new_n1037), .B2(new_n713), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n861), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n788), .A2(new_n370), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n656), .B(new_n1041), .C1(new_n689), .C2(new_n691), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n855), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n861), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n880), .B1(new_n865), .B2(new_n869), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n870), .A2(new_n871), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT104), .B1(new_n877), .B2(KEYINPUT39), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT39), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n874), .B(new_n1049), .C1(new_n876), .C2(new_n865), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1047), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n862), .A2(KEYINPUT116), .A3(new_n881), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT116), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n892), .B1(new_n792), .B2(new_n855), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n880), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1040), .B(new_n1046), .C1(new_n1051), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1046), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT116), .B1(new_n862), .B2(new_n881), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1054), .A2(new_n1053), .A3(new_n880), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1058), .B1(new_n879), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1034), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n861), .B(new_n1063), .C1(new_n712), .C2(new_n887), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1057), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n884), .B1(G330), .B2(new_n896), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n892), .B1(new_n890), .B2(new_n1034), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1068), .A2(new_n1039), .A3(new_n855), .A4(new_n1042), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n856), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1063), .B1(new_n712), .B2(new_n714), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n892), .ZN(new_n1072));
  AOI211_X1 g0872(.A(KEYINPUT117), .B(new_n1070), .C1(new_n1072), .C2(new_n1064), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT117), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1064), .B1(new_n1038), .B2(new_n861), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n856), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1069), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1066), .A2(new_n1067), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1046), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1064), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n1081), .A3(new_n1057), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n674), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT121), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1066), .A2(new_n944), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT118), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1066), .A2(new_n1087), .A3(new_n944), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n738), .A2(new_n202), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n273), .B1(new_n961), .B2(new_n758), .C1(new_n776), .C2(new_n761), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1091), .C1(new_n805), .C2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n753), .A2(G132), .B1(G128), .B2(new_n747), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT119), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n773), .A2(G125), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n736), .A2(new_n813), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n737), .B(new_n1011), .C1(G283), .C2(new_n747), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n266), .B1(new_n760), .B2(new_n777), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n809), .C1(G116), .C2(new_n753), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n756), .A2(new_n210), .B1(new_n212), .B2(new_n758), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1107), .A2(new_n731), .B1(new_n301), .B2(new_n796), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n720), .B(new_n1108), .C1(new_n1051), .C2(new_n729), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1084), .B1(new_n1089), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n944), .ZN(new_n1111));
  AOI211_X1 g0911(.A(KEYINPUT118), .B(new_n1111), .C1(new_n1080), .C2(new_n1057), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1087), .B1(new_n1066), .B2(new_n944), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1084), .B(new_n1109), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1083), .B1(new_n1110), .B2(new_n1115), .ZN(G378));
  INV_X1    g0916(.A(KEYINPUT57), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n889), .A2(G330), .A3(new_n894), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT56), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n320), .A2(new_n310), .A3(new_n829), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT55), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n310), .A2(new_n829), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n313), .A2(new_n316), .A3(new_n319), .A4(new_n1122), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1119), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT55), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(KEYINPUT56), .A3(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1118), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(G330), .A3(new_n889), .A4(new_n894), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n882), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n863), .B1(new_n1051), .B2(new_n880), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1137), .A2(new_n823), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1067), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1066), .B2(new_n1077), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1117), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1081), .B1(new_n1080), .B2(new_n1057), .ZN(new_n1144));
  OAI211_X1 g0944(.A(KEYINPUT57), .B(new_n1143), .C1(new_n1144), .C2(new_n1140), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n674), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1131), .A2(new_n728), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n796), .A2(new_n202), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n801), .A2(new_n1092), .B1(G150), .B2(new_n743), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n754), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n756), .A2(new_n961), .B1(new_n817), .B2(new_n758), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT122), .Z(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(G125), .C2(new_n747), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G41), .B1(new_n803), .B2(G159), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G33), .B1(new_n773), .B2(G124), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n202), .B1(new_n264), .B2(G41), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G116), .A2(new_n747), .B1(new_n769), .B2(G97), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n958), .C1(new_n215), .C2(new_n738), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n736), .A2(new_n207), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n266), .B1(new_n760), .B2(new_n779), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1161), .A2(G41), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n212), .B2(new_n754), .C1(new_n357), .C2(new_n756), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT58), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1158), .A2(new_n1159), .A3(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(new_n731), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT123), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1148), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1169), .B2(new_n1168), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1147), .A2(new_n720), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1143), .B2(new_n944), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1146), .A2(new_n1173), .ZN(G375));
  OR2_X1    g0974(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n925), .A3(new_n1081), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n892), .A2(new_n728), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n756), .A2(new_n212), .B1(new_n224), .B2(new_n758), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT124), .Z(new_n1179));
  AOI22_X1  g0979(.A1(new_n747), .A2(G294), .B1(new_n743), .B2(new_n356), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n273), .B1(new_n773), .B2(G303), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n957), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G283), .B2(new_n753), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1179), .B(new_n1183), .C1(new_n210), .C2(new_n736), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n950), .A2(new_n817), .B1(new_n776), .B2(new_n202), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n266), .B(new_n1185), .C1(new_n769), .C2(new_n1092), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G150), .A2(new_n805), .B1(new_n753), .B2(G137), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G58), .A2(new_n803), .B1(new_n801), .B2(G159), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n760), .A2(new_n1150), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(new_n731), .B1(new_n222), .B2(new_n796), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1177), .A2(new_n720), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1077), .B2(new_n944), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1176), .A2(new_n1194), .ZN(G381));
  NAND3_X1  g0995(.A1(new_n1089), .A2(new_n1083), .A3(new_n1109), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(G375), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G390), .ZN(new_n1199));
  INV_X1    g0999(.A(G384), .ZN(new_n1200));
  INV_X1    g1000(.A(G396), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1003), .A2(new_n1201), .A3(new_n1004), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  OR4_X1    g1004(.A1(G387), .A2(new_n1198), .A3(G381), .A4(new_n1204), .ZN(G407));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1198), .ZN(G409));
  AOI21_X1  g1006(.A(new_n1201), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT125), .B1(new_n1203), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1207), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT125), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1202), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G390), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(G387), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1208), .A2(new_n1211), .A3(G390), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1215), .ZN(new_n1217));
  OAI21_X1  g1017(.A(G387), .B1(new_n1217), .B2(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT62), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT126), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n925), .B(new_n1143), .C1(new_n1144), .C2(new_n1140), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1222), .A2(new_n1173), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n1196), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1173), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1143), .B1(new_n1144), .B2(new_n1140), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n675), .B1(new_n1226), .B2(new_n1117), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1225), .B1(new_n1227), .B2(new_n1145), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1224), .B1(G378), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1221), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1222), .A2(new_n1173), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1233), .A2(new_n1083), .A3(new_n1109), .A4(new_n1089), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1083), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT121), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1237), .B2(new_n1114), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1238), .B2(G375), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1231), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(KEYINPUT126), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1232), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n675), .B1(new_n1175), .B2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1081), .C1(new_n1243), .C2(new_n1175), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(G384), .A3(new_n1194), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G384), .B1(new_n1245), .B2(new_n1194), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1220), .B1(new_n1242), .B2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1239), .A2(new_n1220), .A3(new_n1249), .A4(new_n1240), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1231), .A2(G2897), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1247), .A2(new_n1248), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1232), .A2(new_n1241), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1219), .B1(new_n1250), .B2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1242), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1239), .A2(new_n1249), .A3(new_n1240), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1255), .A2(new_n1256), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1261), .A2(new_n1262), .A3(new_n1252), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1260), .A2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1228), .A2(new_n1196), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(G378), .B2(new_n1228), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1271), .B2(new_n1269), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(new_n1219), .ZN(G402));
endmodule


