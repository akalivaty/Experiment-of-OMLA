//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT66), .B(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT67), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n209), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  AND2_X1   g0023(.A1(KEYINPUT65), .A2(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(KEYINPUT65), .A2(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT64), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n230), .A2(G1), .A3(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n223), .B1(KEYINPUT1), .B2(new_n218), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n220), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G68), .ZN(new_n251));
  INV_X1    g0051(.A(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n250), .B(new_n256), .Z(G351));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G274), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(G226), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n258), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT70), .B(G1698), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(G222), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n229), .A2(new_n231), .B1(G33), .B2(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G77), .B2(new_n273), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n269), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G179), .B2(new_n281), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G150), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n203), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n226), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT71), .A2(G58), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT8), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n229), .A2(new_n231), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n292), .A2(new_n294), .B1(new_n202), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n265), .A2(G20), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n229), .A2(new_n231), .A3(new_n295), .A4(new_n293), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n301));
  OAI211_X1 g0101(.A(G50), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n284), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n281), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n281), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n297), .A2(new_n302), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n297), .B2(new_n302), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT75), .B1(new_n318), .B2(KEYINPUT9), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(KEYINPUT9), .A3(new_n312), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n315), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT10), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n320), .B(new_n321), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n315), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n306), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n291), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n296), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n273), .A2(G226), .A3(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G87), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G1698), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n336), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n334), .B(new_n335), .C1(new_n274), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n279), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n263), .B1(new_n267), .B2(new_n238), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n308), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n342), .B2(new_n279), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(G200), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT79), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n339), .A2(new_n340), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n226), .A2(new_n351), .A3(KEYINPUT7), .ZN(new_n352));
  INV_X1    g0152(.A(G20), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n271), .A2(new_n353), .A3(new_n272), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n252), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n358), .B2(new_n201), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n285), .A2(G159), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n350), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT7), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT78), .B1(new_n339), .B2(new_n340), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT78), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n271), .A2(new_n365), .A3(new_n272), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n252), .B1(new_n354), .B2(KEYINPUT7), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n361), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n371));
  AND4_X1   g0171(.A1(new_n349), .A2(new_n362), .A3(new_n294), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n294), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(KEYINPUT16), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n349), .B1(new_n375), .B2(new_n362), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n333), .B(new_n348), .C1(new_n372), .C2(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n298), .A2(G77), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n299), .A2(new_n379), .B1(G77), .B2(new_n295), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT8), .B(G58), .Z(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n285), .ZN(new_n383));
  INV_X1    g0183(.A(new_n288), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT15), .B(G87), .Z(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(G77), .B2(new_n227), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n380), .B1(new_n387), .B2(new_n294), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n275), .B1(new_n271), .B2(new_n272), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G238), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n390), .B1(new_n206), .B2(new_n273), .C1(new_n238), .C2(new_n341), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n279), .ZN(new_n392));
  INV_X1    g0192(.A(new_n210), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n264), .B1(new_n393), .B2(new_n268), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n388), .B1(new_n282), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(G200), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(new_n388), .C1(new_n308), .C2(new_n395), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n371), .A2(new_n294), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n352), .A2(new_n356), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n406), .B2(new_n370), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT79), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n375), .A2(new_n349), .A3(new_n362), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n332), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n347), .A2(new_n282), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(G179), .B2(new_n347), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n403), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n333), .B1(new_n372), .B2(new_n376), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n347), .A2(G179), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n282), .B2(new_n347), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(KEYINPUT18), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n378), .A2(new_n402), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n252), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n288), .B2(new_n211), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n294), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT11), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n296), .A2(KEYINPUT77), .A3(new_n252), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT12), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT77), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n295), .B2(G68), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n427), .ZN(new_n429));
  INV_X1    g0229(.A(new_n299), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n252), .B1(new_n265), .B2(G20), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n428), .A2(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n336), .A2(new_n338), .A3(G226), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G232), .A2(G1698), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n351), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G97), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n279), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT76), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(KEYINPUT76), .B(new_n279), .C1(new_n438), .C2(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G238), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n263), .B1(new_n267), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n435), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(KEYINPUT13), .B(new_n447), .C1(new_n443), .C2(new_n444), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n434), .B(G169), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n277), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n439), .B1(new_n452), .B2(new_n351), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT76), .B1(new_n453), .B2(new_n279), .ZN(new_n454));
  INV_X1    g0254(.A(new_n444), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n448), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT13), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(new_n435), .A3(new_n448), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(G179), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n458), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n434), .B1(new_n461), .B2(G169), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n433), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G200), .B1(new_n449), .B2(new_n450), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(G190), .A3(new_n458), .ZN(new_n465));
  INV_X1    g0265(.A(new_n433), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n328), .A2(new_n419), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G41), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n265), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(G41), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(KEYINPUT81), .A3(new_n265), .A4(G45), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n476), .ZN(new_n481));
  INV_X1    g0281(.A(new_n474), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n481), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n472), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(G257), .A2(new_n480), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g0287(.A(G244), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n341), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n389), .B2(G250), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT4), .A4(G244), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n279), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(new_n495), .A3(G190), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n486), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G200), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n295), .A2(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n258), .A2(G1), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n299), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(G97), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n206), .B1(new_n352), .B2(new_n356), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n285), .A2(G77), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT80), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  AND4_X1   g0311(.A1(G97), .A2(new_n509), .A3(new_n511), .A4(new_n206), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n509), .A2(new_n511), .B1(new_n207), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n227), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n506), .A2(new_n507), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n504), .B1(new_n516), .B2(new_n294), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n486), .A2(new_n495), .A3(new_n518), .A4(G190), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n497), .A2(new_n499), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n279), .ZN(new_n521));
  OAI211_X1 g0321(.A(G250), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n490), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n341), .A2(new_n488), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(KEYINPUT4), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n525), .B2(new_n489), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n485), .A2(new_n477), .A3(new_n479), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n481), .A2(new_n479), .A3(new_n482), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n260), .ZN(new_n529));
  INV_X1    g0329(.A(G257), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n282), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n509), .A2(new_n511), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n207), .A2(new_n513), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n509), .A2(new_n511), .A3(G97), .A4(new_n206), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n226), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n507), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n505), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n503), .B1(new_n539), .B2(new_n373), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n486), .A2(new_n495), .A3(new_n397), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n532), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n520), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  INV_X1    g0345(.A(G250), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n545), .C1(new_n341), .C2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n480), .A2(G264), .B1(new_n547), .B2(new_n279), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(new_n397), .A3(new_n527), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n279), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n528), .A2(G264), .A3(new_n260), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n527), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n282), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n265), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT25), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT86), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n557), .B(new_n558), .ZN(new_n559));
  OR3_X1    g0359(.A1(new_n555), .A2(KEYINPUT85), .A3(new_n556), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT85), .B1(new_n555), .B2(new_n556), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n299), .A2(new_n501), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n559), .A2(new_n562), .B1(new_n563), .B2(new_n206), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(KEYINPUT65), .A2(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(KEYINPUT65), .A2(G20), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n568), .C1(new_n339), .C2(new_n340), .ZN(new_n569));
  INV_X1    g0369(.A(G87), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n206), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n567), .B2(new_n568), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n575), .A2(G20), .B1(new_n572), .B2(new_n206), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n226), .A2(new_n273), .A3(new_n565), .A4(G87), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n373), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n571), .A2(new_n577), .A3(KEYINPUT24), .A4(new_n578), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n564), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n554), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n502), .A2(G116), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n295), .A2(G116), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n353), .A2(G116), .ZN(new_n588));
  INV_X1    g0388(.A(G283), .ZN(new_n589));
  MUX2_X1   g0389(.A(new_n205), .B(new_n589), .S(G33), .Z(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(new_n226), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n591), .B2(new_n294), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n258), .A2(G97), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n567), .A2(new_n593), .A3(new_n568), .A4(new_n490), .ZN(new_n594));
  INV_X1    g0394(.A(new_n588), .ZN(new_n595));
  AND4_X1   g0395(.A1(KEYINPUT20), .A2(new_n294), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n585), .B(new_n587), .C1(new_n592), .C2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G264), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n271), .A2(G303), .A3(new_n272), .ZN(new_n599));
  OAI21_X1  g0399(.A(G257), .B1(new_n339), .B2(new_n340), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n336), .A2(new_n338), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n279), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n528), .A2(G270), .A3(new_n260), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n527), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n597), .A2(KEYINPUT21), .A3(G169), .A4(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n603), .A2(new_n604), .A3(new_n527), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n597), .A2(new_n607), .A3(G179), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(G270), .A2(new_n480), .B1(new_n483), .B2(new_n485), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n282), .B1(new_n610), .B2(new_n603), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT21), .B1(new_n611), .B2(new_n597), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n584), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n548), .A2(new_n308), .A3(new_n527), .ZN(new_n614));
  INV_X1    g0414(.A(G200), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n552), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n583), .ZN(new_n618));
  NAND2_X1  g0418(.A1(G33), .A2(G116), .ZN(new_n619));
  OAI211_X1 g0419(.A(G244), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n341), .C2(new_n446), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n279), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n265), .A2(new_n484), .A3(G45), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n546), .B1(new_n261), .B2(G1), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n260), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(G169), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g0427(.A(G179), .B(new_n625), .C1(new_n621), .C2(new_n279), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n567), .A2(new_n568), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT83), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n226), .A2(KEYINPUT83), .A3(new_n630), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n570), .A2(new_n205), .A3(new_n206), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n567), .A2(G33), .A3(G97), .A4(new_n568), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT19), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n273), .A2(new_n226), .A3(G68), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n294), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n502), .A2(new_n385), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n385), .A2(new_n295), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n299), .A2(new_n570), .A3(new_n501), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n640), .A3(new_n639), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n644), .B(new_n648), .C1(new_n650), .C2(new_n294), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n625), .B1(new_n621), .B2(new_n279), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n308), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(G200), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n618), .A2(new_n647), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n597), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n308), .B2(new_n605), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n607), .A2(new_n615), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n543), .A2(new_n613), .A3(new_n656), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n471), .A2(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n399), .ZN(new_n664));
  OAI21_X1  g0464(.A(G169), .B1(new_n449), .B2(new_n450), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT14), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n459), .A3(new_n451), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n468), .A2(new_n664), .B1(new_n667), .B2(new_n433), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT17), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n377), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n348), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n418), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n326), .A2(new_n325), .A3(new_n315), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n305), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n515), .A2(new_n507), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n294), .B1(new_n678), .B2(new_n505), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n498), .A2(new_n282), .B1(new_n679), .B2(new_n503), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(new_n655), .A3(new_n647), .A4(new_n541), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .B1(new_n646), .B2(new_n629), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n542), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n651), .A2(new_n654), .B1(new_n629), .B2(new_n646), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n532), .A2(new_n540), .A3(KEYINPUT88), .A4(new_n541), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT87), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n656), .A2(new_n690), .A3(new_n542), .A4(new_n520), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n520), .A2(new_n686), .A3(new_n542), .A4(new_n618), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n613), .B1(new_n692), .B2(KEYINPUT87), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n677), .B1(new_n471), .B2(new_n694), .ZN(G369));
  NOR2_X1   g0495(.A1(new_n609), .A2(new_n612), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n226), .A2(new_n265), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n657), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n696), .B1(new_n660), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n696), .B2(new_n704), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n706), .A2(KEYINPUT89), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(KEYINPUT89), .ZN(new_n708));
  OAI21_X1  g0508(.A(G330), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n579), .A2(new_n580), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n294), .A3(new_n582), .ZN(new_n712));
  INV_X1    g0512(.A(new_n564), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n553), .A3(new_n549), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n702), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n618), .B1(new_n583), .B2(new_n703), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n710), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n696), .A2(new_n702), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n221), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n635), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n234), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n694), .A2(KEYINPUT29), .A3(new_n702), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n486), .A2(new_n495), .A3(new_n548), .A4(new_n652), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n607), .A2(G179), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n526), .A2(new_n531), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n548), .A2(new_n652), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n605), .A2(new_n397), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(KEYINPUT30), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n652), .A2(G179), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n498), .A2(new_n605), .A3(new_n552), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n735), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n742), .A2(new_n743), .A3(new_n702), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n743), .B1(new_n742), .B2(new_n702), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n662), .A2(new_n702), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n684), .A2(KEYINPUT26), .A3(new_n686), .A4(new_n687), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n681), .A2(new_n685), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n647), .B1(new_n692), .B2(new_n613), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n703), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n753), .A2(KEYINPUT29), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n731), .A2(new_n748), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n730), .B1(new_n755), .B2(G1), .ZN(G364));
  AND2_X1   g0556(.A1(new_n226), .A2(G13), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n265), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n724), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n710), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n707), .A2(new_n708), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(G330), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n615), .A2(G190), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n227), .A2(new_n397), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n206), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G58), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n226), .A2(new_n397), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n308), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n767), .B1(new_n768), .B2(new_n771), .C1(new_n211), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n227), .A2(new_n397), .A3(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n775), .A2(KEYINPUT32), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT32), .ZN(new_n778));
  INV_X1    g0578(.A(new_n775), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n779), .B2(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n308), .A2(new_n615), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(G20), .A3(new_n397), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n769), .A2(new_n781), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n273), .B1(new_n570), .B2(new_n782), .C1(new_n783), .C2(new_n202), .ZN(new_n784));
  OR4_X1    g0584(.A1(new_n774), .A2(new_n777), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n226), .B1(new_n397), .B2(new_n770), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n205), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n769), .A2(new_n764), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G68), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  INV_X1    g0591(.A(new_n771), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G322), .A2(new_n792), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n783), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n782), .B(KEYINPUT96), .ZN(new_n797));
  INV_X1    g0597(.A(new_n773), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G303), .A2(new_n797), .B1(new_n798), .B2(G311), .ZN(new_n799));
  INV_X1    g0599(.A(new_n765), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G283), .A2(new_n800), .B1(new_n779), .B2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(new_n786), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n273), .B1(new_n802), .B2(G294), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n785), .A2(new_n791), .B1(new_n796), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n232), .B1(new_n353), .B2(G169), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n256), .A2(new_n261), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT92), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n814), .A2(new_n815), .B1(G45), .B2(new_n234), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n364), .A2(new_n366), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n221), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n816), .B(new_n821), .C1(new_n815), .C2(new_n814), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n273), .A2(new_n221), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G355), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G116), .B2(new_n221), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n813), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n809), .A2(new_n827), .A3(new_n760), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT97), .Z(new_n829));
  INV_X1    g0629(.A(new_n812), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n762), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n763), .A2(new_n831), .ZN(G396));
  NOR2_X1   g0632(.A1(new_n399), .A2(new_n702), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n401), .B1(new_n388), .B2(new_n703), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n399), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n694), .B2(new_n702), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n692), .A2(KEYINPUT87), .ZN(new_n839));
  INV_X1    g0639(.A(new_n613), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n691), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n682), .A2(new_n688), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n402), .A2(new_n703), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n760), .B1(new_n847), .B2(new_n747), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n747), .B2(new_n847), .ZN(new_n849));
  INV_X1    g0649(.A(new_n760), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n808), .A2(new_n810), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n211), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n817), .B1(new_n786), .B2(new_n768), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n797), .A2(G50), .B1(new_n800), .B2(G68), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n775), .ZN(new_n856));
  INV_X1    g0656(.A(new_n783), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G137), .B1(new_n792), .B2(G143), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n788), .C1(new_n776), .C2(new_n773), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n853), .B(new_n856), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n765), .A2(new_n570), .ZN(new_n864));
  INV_X1    g0664(.A(G116), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n773), .A2(new_n865), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(G107), .C2(new_n797), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G294), .A2(new_n792), .B1(new_n779), .B2(G311), .ZN(new_n868));
  INV_X1    g0668(.A(G303), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n868), .B1(new_n589), .B2(new_n788), .C1(new_n869), .C2(new_n783), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n870), .A2(new_n273), .A3(new_n787), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n862), .A2(new_n863), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n837), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n852), .B1(new_n807), .B2(new_n872), .C1(new_n873), .C2(new_n811), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n849), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  NAND2_X1  g0676(.A1(new_n535), .A2(new_n536), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n865), .B(new_n233), .C1(new_n877), .C2(KEYINPUT35), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT35), .B2(new_n877), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OR3_X1    g0680(.A1(new_n234), .A2(new_n358), .A3(new_n211), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n265), .B(G13), .C1(new_n881), .C2(new_n251), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n833), .B1(new_n843), .B2(new_n845), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n433), .A2(new_n702), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n463), .A2(new_n468), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n433), .B(new_n702), .C1(new_n667), .C2(new_n467), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n375), .B1(KEYINPUT16), .B2(new_n374), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n700), .B1(new_n891), .B2(new_n333), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n378), .B2(new_n418), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n333), .ZN(new_n896));
  INV_X1    g0696(.A(new_n700), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n416), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n898), .B2(new_n377), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n408), .A2(new_n409), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n333), .A2(new_n900), .B1(new_n412), .B2(new_n700), .ZN(new_n901));
  INV_X1    g0701(.A(new_n377), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n899), .B1(new_n903), .B2(new_n895), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n894), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n410), .A2(new_n403), .A3(new_n412), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT18), .B1(new_n414), .B2(new_n416), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n892), .B1(new_n909), .B2(new_n672), .ZN(new_n910));
  INV_X1    g0710(.A(new_n899), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n414), .B1(new_n416), .B2(new_n897), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n895), .A3(new_n377), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n906), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n890), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n909), .A2(new_n700), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n667), .A2(new_n433), .A3(new_n703), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT98), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n670), .B(new_n671), .C1(new_n907), .C2(new_n908), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n410), .A2(new_n700), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT99), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n912), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n903), .A2(new_n926), .A3(KEYINPUT37), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT37), .B1(new_n901), .B2(KEYINPUT99), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n902), .B2(new_n901), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n905), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n922), .A2(new_n892), .B1(new_n911), .B2(new_n913), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT39), .B1(new_n932), .B2(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT39), .B1(new_n906), .B2(new_n915), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n921), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n919), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n470), .B1(new_n731), .B2(new_n754), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n677), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n837), .B1(new_n886), .B2(new_n887), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n746), .B(new_n941), .C1(new_n906), .C2(new_n915), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT40), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n941), .A2(KEYINPUT40), .A3(new_n746), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n932), .A2(KEYINPUT38), .ZN(new_n946));
  INV_X1    g0746(.A(new_n923), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n378), .B2(new_n418), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n926), .A2(KEYINPUT37), .B1(new_n377), .B2(new_n912), .ZN(new_n949));
  NOR4_X1   g0749(.A1(new_n901), .A2(new_n902), .A3(new_n925), .A4(new_n895), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n946), .B1(new_n951), .B2(KEYINPUT38), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n470), .A2(new_n746), .ZN(new_n955));
  OAI21_X1  g0755(.A(G330), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n940), .A2(new_n957), .B1(new_n265), .B2(new_n757), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n940), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n883), .B1(new_n958), .B2(new_n959), .ZN(G367));
  INV_X1    g0760(.A(new_n755), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n543), .B1(new_n517), .B2(new_n703), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n680), .A2(new_n541), .A3(new_n702), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n718), .A2(new_n720), .ZN(new_n967));
  INV_X1    g0767(.A(new_n716), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n962), .A2(new_n963), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT44), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT100), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n965), .A2(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n972), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT44), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(KEYINPUT100), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n719), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n719), .B1(new_n974), .B2(new_n977), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n718), .A2(new_n720), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n967), .A2(KEYINPUT101), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n762), .A2(G330), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n709), .A2(KEYINPUT101), .A3(new_n967), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n983), .A3(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n961), .B1(new_n982), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n724), .B(KEYINPUT41), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n758), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n962), .A2(new_n715), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n702), .B1(new_n994), .B2(new_n542), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n964), .A2(new_n718), .A3(new_n720), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(KEYINPUT42), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n686), .B1(new_n651), .B2(new_n703), .ZN(new_n999));
  OR3_X1    g0799(.A1(new_n647), .A2(new_n651), .A3(new_n703), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n997), .A2(new_n998), .B1(KEYINPUT43), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n719), .A2(new_n970), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n993), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n385), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n813), .B1(new_n221), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n820), .A2(new_n244), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n760), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n765), .A2(new_n205), .ZN(new_n1012));
  INV_X1    g0812(.A(G294), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n788), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(G283), .C2(new_n798), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n782), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT46), .B1(new_n1016), .B2(G116), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n817), .B(new_n1017), .C1(G303), .C2(new_n792), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n779), .A2(G317), .B1(new_n802), .B2(G107), .ZN(new_n1019));
  AND2_X1   g0819(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n797), .A2(new_n1020), .B1(new_n857), .B2(G311), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G150), .A2(new_n792), .B1(new_n789), .B2(G159), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G50), .A2(new_n798), .B1(new_n779), .B2(G137), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G143), .A2(new_n857), .B1(new_n800), .B2(G77), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n273), .B1(new_n782), .B2(new_n768), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n802), .B2(G68), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1022), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n807), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1011), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n999), .A2(new_n812), .A3(new_n1000), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1007), .A2(new_n1035), .ZN(G387));
  INV_X1    g0836(.A(new_n989), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n755), .B1(new_n1037), .B2(new_n987), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n988), .A2(new_n961), .A3(new_n989), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n724), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n241), .A2(G45), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT103), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n382), .A2(new_n202), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n726), .B(new_n261), .C1(new_n252), .C2(new_n211), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1042), .B(new_n820), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n824), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(G107), .B2(new_n221), .C1(new_n726), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n850), .B1(new_n1048), .B2(new_n813), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n802), .A2(new_n385), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n771), .B2(new_n202), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT105), .Z(new_n1052));
  AOI211_X1 g0852(.A(new_n818), .B(new_n1012), .C1(G77), .C2(new_n1016), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT104), .B(G150), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n798), .A2(G68), .B1(new_n779), .B2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n857), .A2(G159), .B1(new_n789), .B2(new_n329), .ZN(new_n1056));
  AND4_X1   g0856(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n765), .A2(new_n865), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n818), .B1(new_n775), .B2(new_n795), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n857), .A2(G322), .B1(new_n792), .B2(G317), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n798), .A2(G303), .B1(new_n789), .B2(G311), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT48), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n786), .A2(new_n589), .B1(new_n1013), .B2(new_n782), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT106), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1058), .B(new_n1059), .C1(new_n1067), .C2(KEYINPUT49), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1057), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1049), .B1(new_n1070), .B2(new_n807), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n718), .A2(new_n830), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n990), .B2(new_n759), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1040), .A2(new_n1074), .ZN(G393));
  NOR2_X1   g0875(.A1(new_n964), .A2(new_n830), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT107), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n779), .A2(G322), .B1(G283), .B2(new_n1016), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT108), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n1013), .A2(new_n773), .B1(new_n788), .B2(new_n869), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G116), .B2(new_n802), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1079), .A2(new_n351), .A3(new_n767), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n857), .A2(G317), .B1(new_n792), .B2(G311), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n859), .A2(new_n783), .B1(new_n771), .B2(new_n776), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  AOI211_X1 g0886(.A(new_n818), .B(new_n864), .C1(G68), .C2(new_n1016), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n382), .A2(new_n798), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n802), .A2(G77), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G50), .A2(new_n789), .B1(new_n779), .B2(G143), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1082), .A2(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n808), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n812), .B(new_n808), .C1(G97), .C2(new_n723), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n820), .A2(new_n250), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n850), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1077), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n982), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n724), .B1(new_n1098), .B2(new_n1038), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n982), .B1(new_n755), .B2(new_n990), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1097), .B1(new_n758), .B2(new_n1098), .C1(new_n1099), .C2(new_n1100), .ZN(G390));
  NAND2_X1  g0901(.A1(new_n748), .A2(new_n941), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n921), .B1(new_n884), .B2(new_n889), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n935), .A3(new_n934), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT109), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n888), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n703), .B(new_n836), .C1(new_n751), .C2(new_n752), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n834), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n952), .A3(new_n921), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1105), .A2(KEYINPUT110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT110), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1103), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n934), .A2(new_n935), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT98), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n920), .B(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n834), .B1(new_n694), .B2(new_n844), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n888), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1112), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT110), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1103), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1115), .A2(new_n1124), .A3(new_n759), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT112), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT112), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1115), .A2(new_n1124), .A3(new_n1127), .A4(new_n759), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n938), .B(new_n677), .C1(new_n471), .C2(new_n747), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n873), .A2(new_n746), .A3(G330), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n889), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT111), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n889), .A3(KEYINPUT111), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1102), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1119), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1131), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1109), .B1(new_n748), .B2(new_n941), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1130), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1105), .A2(KEYINPUT110), .A3(new_n1112), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1102), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1146), .B2(new_n1123), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1115), .A2(new_n1124), .A3(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n724), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1116), .A2(new_n811), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n851), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1016), .A2(new_n1054), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G125), .B2(new_n779), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1155), .A2(new_n783), .B1(new_n773), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G137), .B2(new_n789), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n351), .B1(new_n802), .B2(G159), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n792), .A2(G132), .B1(new_n800), .B2(G50), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n773), .A2(new_n205), .B1(new_n775), .B2(new_n1013), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G283), .B2(new_n857), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n273), .B1(new_n800), .B2(G68), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n789), .A2(G107), .B1(new_n802), .B2(G77), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n797), .A2(G87), .B1(new_n792), .B2(G116), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n760), .B1(new_n329), .B2(new_n1151), .C1(new_n1168), .C2(new_n807), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1150), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1129), .A2(new_n1149), .A3(new_n1171), .ZN(G378));
  OAI21_X1  g0972(.A(KEYINPUT115), .B1(new_n919), .B2(new_n936), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n318), .A2(new_n700), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n676), .B2(new_n306), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n305), .B(new_n1176), .C1(new_n674), .C2(new_n675), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n328), .A2(new_n1176), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n676), .A2(new_n306), .A3(new_n1177), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n1174), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n943), .A2(new_n942), .B1(new_n945), .B2(new_n952), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(G330), .ZN(new_n1186));
  AND4_X1   g0986(.A1(G330), .A2(new_n944), .A3(new_n1184), .A4(new_n953), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1173), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1184), .ZN(new_n1189));
  INV_X1    g0989(.A(G330), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n954), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT115), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n890), .A2(new_n916), .B1(new_n909), .B2(new_n700), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1185), .A2(G330), .A3(new_n1184), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1191), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1188), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1130), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1148), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT116), .B1(new_n1200), .B2(KEYINPUT57), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT116), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1123), .B1(new_n1204), .B2(new_n1103), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1130), .B1(new_n1205), .B2(new_n1142), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1202), .B(new_n1203), .C1(new_n1206), .C2(new_n1198), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n937), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1191), .A2(new_n937), .A3(new_n1196), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1203), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1148), .A2(new_n1199), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n725), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1201), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1198), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1189), .A2(new_n810), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n760), .B1(new_n1151), .B2(G50), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G125), .A2(new_n857), .B1(new_n798), .B2(G137), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n792), .A2(G128), .B1(new_n802), .B2(G150), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n855), .B2(new_n788), .C1(new_n782), .C2(new_n1156), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n800), .C2(G159), .ZN(new_n1224));
  INV_X1    g1024(.A(G124), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n775), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT114), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1222), .A2(new_n1223), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n792), .A2(G107), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT113), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n205), .A2(new_n788), .B1(new_n773), .B2(new_n1008), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n768), .A2(new_n765), .B1(new_n775), .B2(new_n589), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n802), .A2(G68), .B1(new_n1016), .B2(G77), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n818), .A2(new_n259), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G116), .B2(new_n857), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1230), .A2(new_n1233), .A3(new_n1234), .A4(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT58), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1235), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1228), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1217), .B1(new_n1242), .B2(new_n808), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1215), .A2(new_n759), .B1(new_n1216), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1214), .A2(new_n1244), .ZN(G375));
  INV_X1    g1045(.A(new_n992), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1136), .A2(new_n1119), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1130), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1143), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n797), .A2(G97), .B1(new_n792), .B2(G283), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1050), .C1(new_n865), .C2(new_n788), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n273), .B(new_n1251), .C1(G77), .C2(new_n800), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n783), .A2(new_n1013), .B1(new_n775), .B2(new_n869), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G107), .B2(new_n798), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n773), .A2(new_n859), .B1(new_n786), .B2(new_n202), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT117), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n797), .A2(G159), .B1(new_n792), .B2(G137), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1155), .B2(new_n775), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n817), .B1(new_n765), .B2(new_n768), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n855), .A2(new_n783), .B1(new_n788), .B2(new_n1156), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1252), .A2(new_n1254), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n760), .B1(G68), .B2(new_n1151), .C1(new_n1262), .C2(new_n807), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1138), .B2(new_n810), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1247), .B2(new_n758), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1249), .A2(new_n1267), .ZN(G381));
  OR2_X1    g1068(.A1(G390), .A2(G384), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1040), .A2(new_n1074), .A3(new_n831), .A4(new_n763), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1269), .A2(G387), .A3(G381), .A4(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT118), .Z(new_n1272));
  OR3_X1    g1072(.A1(new_n1272), .A2(G378), .A3(G375), .ZN(G407));
  NAND2_X1  g1073(.A1(new_n701), .A2(G213), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(G375), .A2(G378), .A3(new_n1274), .ZN(new_n1275));
  XOR2_X1   g1075(.A(new_n1275), .B(KEYINPUT119), .Z(new_n1276));
  NAND3_X1  g1076(.A1(G407), .A2(G213), .A3(new_n1276), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(new_n1270), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1278), .A3(new_n1270), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n993), .A2(new_n1006), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1281), .B(new_n1282), .C1(new_n1283), .C2(KEYINPUT124), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1282), .ZN(new_n1285));
  OAI21_X1  g1085(.A(G387), .B1(new_n1285), .B2(new_n1280), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1284), .A2(new_n1286), .A3(G390), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G390), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1214), .A2(G378), .A3(new_n1244), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT120), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1186), .A2(new_n1187), .A3(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n759), .B1(new_n1294), .B2(new_n1208), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1216), .A2(new_n1243), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1246), .B2(new_n1200), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1292), .B1(new_n1298), .B2(G378), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1212), .A2(new_n1215), .A3(new_n1246), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1115), .A2(new_n1124), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n725), .B1(new_n1303), .B2(new_n1143), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1170), .B1(new_n1304), .B2(new_n1148), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1302), .A2(KEYINPUT120), .A3(new_n1129), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1299), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1274), .B1(new_n1291), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT60), .B1(new_n1247), .B2(new_n1130), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1248), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1247), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n724), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT121), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n725), .B1(new_n1309), .B2(new_n1248), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT121), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1311), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1317), .B2(new_n1267), .ZN(new_n1318));
  AOI211_X1 g1118(.A(new_n875), .B(new_n1266), .C1(new_n1313), .C2(new_n1316), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n701), .A2(G213), .A3(G2897), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1312), .A2(KEYINPUT121), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1315), .B1(new_n1314), .B2(new_n1311), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1267), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n875), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1317), .A2(G384), .A3(new_n1267), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1320), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1322), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1290), .B1(new_n1308), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1274), .B(new_n1331), .C1(new_n1291), .C2(new_n1307), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(KEYINPUT122), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1330), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1214), .A2(G378), .A3(new_n1244), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1299), .A3(new_n1306), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1338), .A2(KEYINPUT122), .A3(new_n1274), .A4(new_n1331), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT62), .B1(new_n1339), .B2(KEYINPUT126), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1289), .B1(new_n1336), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1342), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1343), .B1(new_n1308), .B2(new_n1329), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT63), .ZN(new_n1345));
  OR2_X1    g1145(.A1(new_n1332), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT122), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1332), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1339), .A2(new_n1345), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1344), .B(new_n1346), .C1(new_n1348), .C2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1341), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT127), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1341), .A2(new_n1350), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(G405));
  XOR2_X1   g1155(.A(G375), .B(G378), .Z(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1331), .ZN(new_n1357));
  XNOR2_X1  g1157(.A(new_n1357), .B(new_n1289), .ZN(G402));
endmodule


