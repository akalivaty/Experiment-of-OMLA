//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  OAI211_X1 g010(.A(G128), .B(new_n193), .C1(new_n194), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(new_n199), .C1(KEYINPUT1), .C2(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n202), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n197), .A2(new_n201), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n213), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT79), .B1(new_n217), .B2(new_n218), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT11), .A3(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n232), .A2(new_n224), .A3(new_n226), .A4(new_n227), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n221), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT12), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n221), .A2(KEYINPUT12), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT77), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n204), .A2(new_n207), .A3(new_n242), .A4(new_n209), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(G101), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n210), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n245), .A3(G101), .A4(new_n243), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n241), .A2(new_n250), .A3(G101), .A4(new_n243), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n198), .A2(new_n199), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n198), .A2(new_n199), .A3(new_n252), .A4(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT0), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n200), .A3(KEYINPUT65), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(KEYINPUT0), .B2(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n252), .B1(new_n198), .B2(new_n199), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n254), .A2(new_n256), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n251), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n249), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n234), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT10), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n216), .A2(new_n268), .A3(new_n220), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n202), .A2(new_n214), .A3(KEYINPUT10), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(new_n267), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n191), .B1(new_n239), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n250), .B1(new_n244), .B2(new_n246), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n264), .B1(new_n274), .B2(new_n248), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n234), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n276), .A2(new_n271), .A3(new_n191), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT80), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n271), .A3(new_n191), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n273), .A2(new_n275), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n267), .A2(new_n281), .B1(new_n237), .B2(new_n238), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n279), .B(new_n280), .C1(new_n282), .C2(new_n191), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(G469), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n239), .A2(new_n191), .A3(new_n271), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n191), .B1(new_n276), .B2(new_n271), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(KEYINPUT81), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT81), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n290), .B(new_n191), .C1(new_n276), .C2(new_n271), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n285), .B(new_n286), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(G469), .A2(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  OAI21_X1  g109(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT76), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G472), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n228), .A2(new_n229), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n225), .A2(G134), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n227), .A3(G131), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(KEYINPUT69), .A3(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n202), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G116), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n263), .A2(new_n319), .A3(new_n234), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n263), .B2(new_n234), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n308), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n263), .A2(new_n234), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n202), .A2(new_n304), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n317), .B1(new_n263), .B2(new_n234), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT28), .B1(new_n308), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G237), .ZN(new_n335));
  AOI21_X1  g149(.A(G953), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G210), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n339), .A3(G210), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G101), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n338), .B2(new_n340), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n328), .A2(new_n331), .A3(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n308), .B(KEYINPUT30), .C1(new_n320), .C2(new_n321), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n347));
  NAND2_X1  g161(.A1(new_n325), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n317), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n322), .ZN(new_n350));
  INV_X1    g164(.A(new_n344), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n308), .B1(new_n320), .B2(new_n321), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n317), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n322), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n330), .B1(new_n357), .B2(KEYINPUT28), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n351), .A2(new_n353), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n300), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT31), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n322), .A2(KEYINPUT71), .A3(new_n344), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT71), .B1(new_n322), .B2(new_n344), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT31), .A3(new_n349), .A4(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n344), .B1(new_n328), .B2(new_n331), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(G472), .A2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n363), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n368), .B2(new_n370), .ZN(new_n377));
  INV_X1    g191(.A(new_n375), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n377), .A2(KEYINPUT32), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n362), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(G234), .B2(new_n286), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n309), .B2(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n385), .B(new_n386), .C1(G119), .C2(new_n200), .ZN(new_n387));
  XNOR2_X1  g201(.A(G119), .B(G128), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT24), .B(G110), .Z(new_n389));
  AOI22_X1  g203(.A1(new_n387), .A2(G110), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G125), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G125), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n394), .A3(G140), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n391), .A2(G140), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT73), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT73), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n400), .A3(KEYINPUT16), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT72), .B(G125), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(KEYINPUT16), .A3(G140), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(G146), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AOI211_X1 g220(.A(new_n195), .B(new_n404), .C1(new_n399), .C2(new_n401), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n390), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(G146), .A3(new_n405), .ZN(new_n409));
  XNOR2_X1  g223(.A(G125), .B(G140), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT74), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n195), .ZN(new_n412));
  OAI22_X1  g226(.A1(new_n387), .A2(G110), .B1(new_n388), .B2(new_n389), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G953), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(G221), .A3(G234), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT75), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT22), .B(G137), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n408), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n408), .B2(new_n414), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n286), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT25), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n408), .A2(new_n414), .ZN(new_n426));
  INV_X1    g240(.A(new_n419), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n420), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT25), .A3(new_n286), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n383), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n382), .A2(G902), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n299), .A2(new_n380), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G224), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G953), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n263), .A2(new_n403), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n217), .A2(new_n403), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI221_X1 g256(.A(new_n440), .B1(new_n437), .B2(G953), .C1(new_n263), .C2(new_n403), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n251), .A2(new_n317), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n274), .B2(new_n248), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT5), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(G113), .C1(KEYINPUT5), .C2(new_n310), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n315), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n218), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n447), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n449), .A2(new_n447), .A3(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n456), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n447), .B(new_n458), .C1(new_n449), .C2(new_n453), .ZN(new_n459));
  AOI211_X1 g273(.A(KEYINPUT83), .B(new_n445), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n461));
  INV_X1    g275(.A(new_n448), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n453), .B1(new_n249), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n456), .B1(new_n463), .B2(new_n446), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n446), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n461), .B1(new_n466), .B2(new_n444), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n451), .A2(new_n315), .B1(new_n210), .B2(new_n213), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n446), .B(KEYINPUT8), .Z(new_n471));
  OAI21_X1  g285(.A(KEYINPUT84), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n452), .A2(new_n218), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n214), .A2(new_n315), .A3(new_n451), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n438), .A2(KEYINPUT7), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n444), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n439), .B2(new_n441), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n478), .A2(new_n481), .A3(new_n486), .A4(new_n482), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n249), .A2(new_n462), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n446), .A3(new_n474), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n286), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n436), .B1(new_n468), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n463), .A2(new_n446), .A3(new_n456), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n458), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n454), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT83), .B1(new_n495), .B2(new_n445), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n466), .A2(new_n461), .A3(new_n444), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n487), .A2(new_n489), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n499), .B2(new_n484), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n500), .A3(new_n435), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n311), .A2(G122), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(KEYINPUT14), .ZN(new_n505));
  INV_X1    g319(.A(G122), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G116), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(KEYINPUT14), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n504), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n510));
  OAI21_X1  g324(.A(G107), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n200), .A2(G143), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n192), .A2(G128), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n223), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n504), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n507), .B2(new_n504), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n206), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n223), .ZN(new_n522));
  INV_X1    g336(.A(new_n519), .ZN(new_n523));
  AOI21_X1  g337(.A(G107), .B1(new_n523), .B2(new_n517), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n518), .A2(new_n206), .A3(new_n519), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n192), .A2(G128), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n529), .A2(KEYINPUT89), .B1(KEYINPUT13), .B2(new_n512), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n527), .C1(new_n513), .C2(new_n528), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n223), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n521), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n295), .A2(new_n381), .A3(G953), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n523), .A2(G107), .A3(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n520), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n530), .A2(new_n532), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n522), .B(new_n539), .C1(new_n540), .C2(new_n223), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n535), .B1(new_n541), .B2(new_n521), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n286), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G478), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n543), .B(new_n545), .Z(new_n546));
  XNOR2_X1  g360(.A(G113), .B(G122), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(new_n203), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n334), .A2(G237), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n550));
  OAI211_X1 g364(.A(G214), .B(new_n415), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n192), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n229), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT86), .ZN(new_n555));
  INV_X1    g369(.A(new_n553), .ZN(new_n556));
  AOI21_X1  g370(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n557));
  OAI21_X1  g371(.A(G131), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n552), .A2(new_n559), .A3(new_n553), .A4(new_n229), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n411), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n396), .B1(new_n403), .B2(G140), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n561), .B(new_n409), .C1(G146), .C2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n412), .B1(new_n195), .B2(new_n564), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT18), .B(G131), .C1(new_n556), .C2(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(KEYINPUT18), .A2(G131), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n552), .A2(new_n553), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n548), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n575), .B(new_n229), .C1(new_n552), .C2(new_n553), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n406), .A2(new_n407), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n555), .A2(new_n575), .A3(new_n558), .A4(new_n560), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT87), .B1(new_n579), .B2(new_n548), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n402), .A2(new_n405), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n195), .ZN(new_n582));
  INV_X1    g396(.A(new_n576), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n578), .A2(new_n582), .A3(new_n409), .A4(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT87), .A3(new_n548), .A4(new_n571), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n573), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT20), .ZN(new_n588));
  NOR2_X1   g402(.A1(G475), .A2(G902), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n548), .A3(new_n571), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n572), .B1(new_n593), .B2(new_n585), .ZN(new_n594));
  INV_X1    g408(.A(new_n589), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT20), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n584), .A2(new_n571), .ZN(new_n597));
  INV_X1    g411(.A(new_n548), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n580), .B2(new_n586), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n286), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n590), .A2(new_n596), .B1(new_n601), .B2(G475), .ZN(new_n602));
  NAND2_X1  g416(.A1(G234), .A2(G237), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(G952), .A3(new_n415), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(G902), .A3(G953), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT21), .B(G898), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G214), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n502), .A2(new_n546), .A3(new_n602), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n434), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n208), .ZN(G3));
  OAI21_X1  g429(.A(G472), .B1(new_n377), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n374), .A2(new_n375), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n299), .A2(new_n619), .A3(KEYINPUT91), .A4(new_n433), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT91), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n294), .A2(new_n298), .A3(new_n617), .A4(new_n616), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT25), .B1(new_n429), .B2(new_n286), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n424), .B(G902), .C1(new_n428), .C2(new_n420), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n382), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n429), .ZN(new_n626));
  INV_X1    g440(.A(new_n432), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n621), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT92), .Z(new_n631));
  INV_X1    g445(.A(new_n609), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n544), .A2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n534), .A2(new_n536), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n541), .A2(new_n521), .A3(new_n535), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n633), .B(new_n634), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n634), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n537), .B2(new_n542), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n638), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT94), .B1(new_n543), .B2(new_n544), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT95), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n641), .B(new_n648), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n602), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n435), .B1(new_n498), .B2(new_n500), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT93), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n611), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n492), .A2(KEYINPUT93), .A3(new_n501), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n631), .A2(new_n632), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n203), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NAND2_X1  g475(.A1(new_n590), .A2(new_n596), .ZN(new_n662));
  INV_X1    g476(.A(new_n546), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n601), .A2(G475), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n654), .A3(new_n655), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n631), .A2(new_n632), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n408), .A2(new_n673), .A3(new_n414), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n673), .B1(new_n408), .B2(new_n414), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n675), .A2(new_n676), .B1(KEYINPUT36), .B2(new_n419), .ZN(new_n677));
  INV_X1    g491(.A(new_n676), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n419), .A2(KEYINPUT36), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n674), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n627), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n672), .B1(new_n431), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n625), .A2(new_n683), .A3(KEYINPUT98), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n299), .A2(new_n619), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n613), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT37), .B(G110), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  OR2_X1    g503(.A1(new_n606), .A2(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n604), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n299), .A2(new_n380), .A3(new_n685), .A4(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n667), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n200), .ZN(G30));
  XNOR2_X1  g508(.A(new_n691), .B(KEYINPUT39), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n294), .A2(new_n298), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT40), .Z(new_n697));
  NAND3_X1  g511(.A1(new_n374), .A2(new_n363), .A3(new_n375), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT32), .B1(new_n377), .B2(new_n378), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n369), .A2(new_n349), .A3(new_n365), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n357), .A2(new_n351), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n700), .B1(new_n300), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n682), .A2(new_n684), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n602), .A2(new_n546), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n610), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n502), .B(KEYINPUT38), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n697), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  NOR2_X1   g524(.A1(new_n692), .A2(new_n656), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n195), .ZN(G48));
  AND2_X1   g526(.A1(new_n654), .A2(new_n655), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n361), .B1(new_n698), .B2(new_n699), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n286), .B1(new_n289), .B2(new_n291), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n296), .A3(new_n292), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n714), .A2(new_n628), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n713), .A2(new_n632), .A3(new_n718), .A4(new_n651), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND3_X1  g535(.A1(new_n668), .A2(new_n632), .A3(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AND3_X1   g537(.A1(new_n716), .A2(new_n296), .A3(new_n292), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n654), .A2(new_n655), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT99), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT99), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n654), .A2(new_n655), .A3(new_n727), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n662), .A2(new_n546), .A3(new_n664), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n380), .A3(new_n632), .A4(new_n685), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT100), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n735), .B(new_n732), .C1(new_n726), .C2(new_n728), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n309), .ZN(G21));
  NAND3_X1  g552(.A1(new_n706), .A2(new_n654), .A3(new_n655), .ZN(new_n739));
  INV_X1    g553(.A(new_n321), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n263), .A2(new_n319), .A3(new_n234), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n318), .B1(new_n742), .B2(new_n308), .ZN(new_n743));
  INV_X1    g557(.A(new_n322), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT28), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n331), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n351), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n371), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n375), .B(KEYINPUT101), .Z(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(KEYINPUT102), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n368), .A2(new_n370), .B1(new_n746), .B2(new_n351), .ZN(new_n752));
  INV_X1    g566(.A(new_n749), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n374), .A2(new_n286), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n750), .A2(new_n754), .B1(new_n755), .B2(G472), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n632), .A3(new_n724), .A4(new_n433), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n739), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n506), .ZN(G24));
  INV_X1    g573(.A(new_n691), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n602), .A2(new_n650), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n685), .A3(new_n756), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n726), .B2(new_n728), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n391), .ZN(G27));
  INV_X1    g578(.A(new_n296), .ZN(new_n765));
  INV_X1    g579(.A(new_n238), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT12), .B1(new_n221), .B2(new_n234), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n271), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n190), .B1(new_n281), .B2(new_n267), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n190), .A2(new_n768), .B1(new_n769), .B2(new_n276), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n770), .B2(G902), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n765), .B1(new_n292), .B2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n492), .A2(new_n772), .A3(new_n501), .A4(new_n610), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n628), .B1(new_n700), .B2(new_n362), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n761), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n774), .A3(new_n761), .A4(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT103), .B(G131), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G33));
  NAND4_X1  g595(.A1(new_n773), .A2(new_n774), .A3(new_n666), .A4(new_n691), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT104), .B(G134), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G36));
  NAND2_X1  g598(.A1(new_n662), .A2(new_n664), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT43), .B1(new_n785), .B2(new_n650), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n647), .A2(new_n649), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n602), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n786), .A2(new_n618), .A3(new_n789), .A4(new_n685), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n695), .ZN(new_n793));
  INV_X1    g607(.A(new_n292), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n770), .A2(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(G469), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT45), .B1(new_n278), .B2(new_n283), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n293), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT46), .B(new_n293), .C1(new_n796), .C2(new_n797), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n765), .B(new_n793), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n705), .A2(new_n619), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT44), .A3(new_n786), .A4(new_n789), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n502), .A2(new_n611), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n792), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  AOI21_X1  g621(.A(new_n765), .B1(new_n800), .B2(new_n801), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n380), .A2(new_n433), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n761), .A3(new_n805), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n692), .B1(new_n656), .B2(new_n667), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n763), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n431), .A2(new_n681), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n292), .A2(new_n771), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n821), .A2(new_n822), .A3(new_n765), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n704), .A2(new_n819), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n739), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n816), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n763), .A2(new_n817), .A3(new_n825), .A4(KEYINPUT52), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n815), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n651), .A2(new_n756), .A3(new_n685), .A4(new_n691), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n729), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n817), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n826), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n818), .A2(new_n816), .A3(new_n826), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT107), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n613), .B1(new_n434), .B2(new_n686), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n758), .ZN(new_n838));
  INV_X1    g652(.A(new_n501), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n612), .B1(new_n839), .B2(new_n652), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n665), .B1(new_n602), .B2(new_n650), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n620), .A2(new_n629), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n838), .A2(new_n719), .A3(new_n722), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n294), .A2(new_n298), .A3(new_n691), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n705), .A2(new_n845), .A3(new_n714), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n502), .A2(new_n730), .A3(new_n611), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n830), .A2(new_n773), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n779), .A2(new_n848), .A3(new_n782), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n737), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n829), .A2(new_n836), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n834), .A4(new_n835), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n829), .A2(new_n836), .A3(new_n850), .A4(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n834), .A2(new_n835), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n779), .A2(new_n782), .A3(new_n848), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n840), .A2(new_n730), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n294), .A2(new_n298), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n714), .A2(new_n861), .A3(new_n628), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n705), .A2(new_n622), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n750), .A2(new_n754), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n433), .A3(new_n616), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n716), .A2(new_n632), .A3(new_n296), .A4(new_n292), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n713), .A3(new_n706), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n719), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n841), .A2(new_n842), .ZN(new_n871));
  INV_X1    g685(.A(new_n718), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n666), .A2(new_n654), .A3(new_n655), .A4(new_n632), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n630), .A2(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n859), .B(new_n875), .C1(new_n734), .C2(new_n736), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n852), .B1(new_n858), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n857), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT109), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT109), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n857), .A2(new_n881), .A3(new_n877), .A4(new_n878), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n786), .A2(new_n605), .A3(new_n789), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n883), .A2(KEYINPUT110), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(KEYINPUT110), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n866), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(KEYINPUT111), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n708), .A2(new_n610), .A3(new_n717), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(KEYINPUT111), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n886), .B(new_n889), .C1(KEYINPUT111), .C2(new_n887), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n704), .A2(new_n604), .A3(new_n628), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n502), .A2(new_n611), .A3(new_n717), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n896), .A2(new_n785), .A3(new_n787), .ZN(new_n897));
  INV_X1    g711(.A(new_n895), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n884), .B2(new_n885), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n756), .A2(new_n685), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n716), .A2(new_n292), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n297), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n809), .A2(new_n810), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n886), .A2(new_n905), .A3(new_n805), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n892), .A2(new_n893), .A3(new_n902), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT51), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n884), .A2(new_n885), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n774), .A3(new_n895), .ZN(new_n911));
  XOR2_X1   g725(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n912));
  OR2_X1    g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  INV_X1    g728(.A(new_n651), .ZN(new_n915));
  OAI211_X1 g729(.A(G952), .B(new_n415), .C1(new_n896), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n886), .B2(new_n729), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n900), .B(new_n898), .C1(new_n884), .C2(new_n885), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT112), .B1(new_n920), .B2(new_n897), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n899), .A2(new_n901), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT112), .ZN(new_n923));
  INV_X1    g737(.A(new_n897), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n921), .A2(new_n925), .A3(new_n892), .A4(new_n893), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT113), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n886), .B(new_n805), .C1(new_n905), .C2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n905), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT51), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n919), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n856), .A2(new_n880), .A3(new_n882), .A4(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(G952), .A2(G953), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n433), .A2(new_n610), .A3(new_n298), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT105), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n704), .ZN(new_n938));
  INV_X1    g752(.A(new_n708), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n785), .A2(new_n650), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n903), .B(KEYINPUT49), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n935), .A2(new_n942), .ZN(G75));
  NOR2_X1   g757(.A1(new_n415), .A2(G952), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n857), .A2(new_n877), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n946), .A2(G210), .A3(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n466), .B(new_n444), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(KEYINPUT56), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n945), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(G210), .A3(G902), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT115), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n286), .B1(new_n857), .B2(new_n877), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(KEYINPUT115), .A3(G210), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n951), .B1(new_n958), .B2(new_n949), .ZN(G51));
  NOR2_X1   g773(.A1(new_n796), .A2(new_n797), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n956), .A2(KEYINPUT116), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT116), .B1(new_n956), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n293), .B(KEYINPUT57), .Z(new_n964));
  AND3_X1   g778(.A1(new_n857), .A2(new_n877), .A3(new_n878), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n878), .B1(new_n857), .B2(new_n877), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n289), .A2(new_n291), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n944), .B1(new_n963), .B2(new_n969), .ZN(G54));
  AND2_X1   g784(.A1(KEYINPUT58), .A2(G475), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n946), .A2(G902), .A3(new_n587), .A4(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT117), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n956), .A2(new_n971), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n944), .B1(new_n976), .B2(new_n594), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(G60));
  NOR2_X1   g792(.A1(new_n639), .A2(new_n640), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  NOR2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n965), .B2(new_n966), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n945), .ZN(new_n984));
  INV_X1    g798(.A(new_n981), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n858), .A2(new_n876), .A3(new_n852), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n852), .B2(new_n851), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT54), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n882), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n879), .A2(KEYINPUT109), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n984), .B1(new_n991), .B2(new_n979), .ZN(G63));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT119), .ZN(new_n995));
  XNOR2_X1  g809(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n857), .B2(new_n877), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n677), .A2(new_n680), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT120), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n945), .B1(new_n999), .B2(new_n429), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n993), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n999), .A2(new_n429), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1006), .A2(KEYINPUT61), .A3(new_n945), .A4(new_n1002), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(G66));
  OAI21_X1  g822(.A(G953), .B1(new_n608), .B2(new_n437), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n875), .B1(new_n734), .B2(new_n736), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1010), .A2(KEYINPUT121), .A3(new_n415), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT121), .B1(new_n1010), .B2(new_n415), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT122), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n495), .B1(G898), .B2(new_n415), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1014), .B(new_n1016), .ZN(G69));
  INV_X1    g831(.A(new_n696), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n805), .A2(new_n842), .A3(new_n774), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT124), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(KEYINPUT125), .A3(new_n806), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(KEYINPUT125), .B1(new_n1021), .B2(new_n806), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n813), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n831), .A2(new_n832), .ZN(new_n1026));
  INV_X1    g840(.A(new_n709), .ZN(new_n1027));
  OAI21_X1  g841(.A(KEYINPUT62), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT62), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n818), .A2(new_n1029), .A3(new_n709), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(KEYINPUT126), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT126), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1035));
  INV_X1    g849(.A(new_n806), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1019), .B(KEYINPUT124), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n1022), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1033), .A2(new_n1034), .A3(new_n813), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n346), .A2(new_n348), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n565), .B(KEYINPUT123), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1041), .A2(new_n415), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n188), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n415), .B1(new_n1046), .B2(G900), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n802), .A2(new_n774), .A3(new_n713), .A4(new_n706), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n813), .A2(new_n806), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n818), .A2(new_n779), .A3(new_n782), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n415), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1044), .B1(new_n188), .B2(G953), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1047), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1045), .A2(new_n1053), .ZN(G72));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  INV_X1    g870(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1010), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n349), .A2(new_n322), .A3(new_n351), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n945), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n350), .A2(new_n344), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n1032), .A2(new_n1040), .A3(new_n1059), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1063), .B1(new_n1064), .B2(new_n1056), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1057), .B1(new_n701), .B2(new_n352), .ZN(new_n1066));
  INV_X1    g880(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g881(.A(KEYINPUT127), .B1(new_n987), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(KEYINPUT127), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n855), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1070));
  AOI211_X1 g884(.A(new_n1062), .B(new_n1065), .C1(new_n1068), .C2(new_n1070), .ZN(G57));
endmodule


