//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n461), .B2(new_n462), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n482), .B(new_n485), .C1(new_n462), .C2(new_n461), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT66), .A2(G114), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT66), .A2(G114), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n488), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(KEYINPUT66), .A2(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT66), .A2(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n465), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT67), .B1(new_n495), .B2(new_n465), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n491), .B(G2104), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n487), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT69), .ZN(new_n504));
  OAI21_X1  g079(.A(G651), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n505), .B1(new_n517), .B2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(new_n513), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n506), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(G51), .B1(new_n501), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n522), .B(new_n530), .C1(new_n523), .C2(new_n513), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n507), .A2(new_n537), .B1(new_n513), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  XOR2_X1   g115(.A(KEYINPUT71), .B(G43), .Z(new_n541));
  INV_X1    g116(.A(new_n513), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n527), .A2(new_n541), .B1(new_n542), .B2(G81), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n535), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT72), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT74), .B1(new_n513), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n507), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n506), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n510), .A2(new_n509), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n558), .A2(new_n563), .A3(new_n568), .ZN(G299));
  OR2_X1    g144(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n527), .A2(G49), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n542), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  OAI21_X1  g150(.A(G61), .B1(new_n510), .B2(new_n509), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(KEYINPUT75), .B(G61), .C1(new_n510), .C2(new_n509), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT76), .B1(new_n513), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n501), .A2(new_n506), .A3(new_n585), .A4(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(G48), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n506), .A2(new_n590), .A3(G48), .A4(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n582), .A2(new_n587), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n535), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n507), .A2(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n595), .B2(new_n598), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n513), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n527), .A2(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  INV_X1    g186(.A(G79), .ZN(new_n612));
  INV_X1    g187(.A(G543), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n565), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI221_X1 g191(.A(KEYINPUT79), .B1(new_n612), .B2(new_n613), .C1(new_n565), .C2(new_n611), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n616), .A2(G651), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n603), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n603), .B1(new_n620), .B2(G868), .ZN(G321));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(G299), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(G168), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(new_n623), .B2(G168), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g207(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n464), .A2(G135), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT80), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n475), .B2(G123), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n635), .A2(new_n636), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n639), .A2(new_n644), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n637), .A2(new_n645), .A3(new_n646), .A4(new_n648), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n636), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n640), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT81), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n678), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n682), .A3(new_n678), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n683), .B1(new_n682), .B2(new_n678), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G6), .A2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G305), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT86), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n703), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G1971), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  NOR2_X1   g287(.A1(new_n706), .A2(G1971), .ZN(new_n713));
  NOR4_X1   g288(.A1(new_n702), .A2(new_n707), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n464), .A2(G131), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  INV_X1    g298(.A(G107), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G2105), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n475), .B2(G119), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n719), .B1(new_n727), .B2(new_n718), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT84), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n703), .A2(G24), .ZN(new_n734));
  INV_X1    g309(.A(G290), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n703), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1986), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n716), .A2(new_n717), .A3(new_n732), .A4(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT36), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT36), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G171), .A2(new_n703), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G5), .B2(new_n703), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT97), .Z(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2078), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G168), .A2(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(KEYINPUT94), .C1(G16), .C2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT94), .B2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT95), .B(G1966), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n547), .A2(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G16), .B2(G19), .ZN(new_n758));
  INV_X1    g333(.A(G1341), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G162), .A2(G29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G29), .B2(G35), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT29), .B(G2090), .Z(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT31), .B(G11), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n718), .B1(new_n768), .B2(G28), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n767), .B1(new_n769), .B2(new_n770), .C1(new_n647), .C2(new_n718), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n758), .B2(new_n759), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n744), .A2(new_n745), .B1(new_n762), .B2(new_n763), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(G34), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n718), .B1(new_n774), .B2(G34), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n472), .A2(new_n718), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2084), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n765), .A2(new_n772), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n475), .A2(G129), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT26), .Z(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n784), .A2(KEYINPUT93), .A3(new_n718), .ZN(new_n785));
  INV_X1    g360(.A(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G29), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G29), .B2(G32), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT27), .B(G1996), .Z(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n703), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1956), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n718), .A2(G26), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT28), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n464), .A2(G140), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n475), .A2(G128), .ZN(new_n800));
  OR2_X1    g375(.A1(G104), .A2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(new_n718), .ZN(new_n805));
  INV_X1    g380(.A(G2067), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n790), .A2(new_n791), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n792), .A2(new_n796), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n751), .A2(new_n756), .A3(new_n779), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G4), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n620), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT88), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT87), .B(G1348), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n718), .A2(G33), .ZN(new_n817));
  NAND2_X1  g392(.A1(G115), .A2(G2104), .ZN(new_n818));
  INV_X1    g393(.A(G127), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n463), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n465), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n824));
  NAND2_X1  g399(.A1(G103), .A2(G2104), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(G2105), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n464), .A2(G139), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n817), .B1(new_n829), .B2(new_n718), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT90), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G2072), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT91), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(G2072), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n742), .A2(new_n816), .A3(new_n837), .ZN(G311));
  NAND3_X1  g413(.A1(new_n742), .A2(new_n816), .A3(new_n837), .ZN(G150));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n565), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g419(.A(KEYINPUT98), .B(new_n840), .C1(new_n565), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(G651), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT99), .B(G93), .ZN(new_n847));
  AOI22_X1  g422(.A1(G55), .A2(new_n527), .B1(new_n542), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n620), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n849), .A2(new_n546), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n846), .A2(new_n543), .A3(new_n848), .A4(new_n545), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n857), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT39), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT39), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(G145));
  NAND2_X1  g441(.A1(new_n464), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n475), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n727), .A2(KEYINPUT102), .ZN(new_n872));
  INV_X1    g447(.A(new_n634), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n722), .A2(new_n726), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n873), .B1(new_n872), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(new_n871), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n499), .B(new_n803), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n784), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n829), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n829), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n472), .B(new_n479), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n647), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n888), .A2(new_n880), .A3(new_n883), .A4(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n886), .A2(new_n829), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(new_n887), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n884), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n893), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n884), .B2(new_n899), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n895), .B(new_n896), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n884), .A2(new_n899), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n890), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n901), .A3(new_n900), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(KEYINPUT104), .A3(new_n896), .A4(new_n895), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT40), .B1(new_n906), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(G395));
  XNOR2_X1  g488(.A(new_n629), .B(new_n857), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n556), .A2(new_n557), .B1(G651), .B2(new_n567), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n563), .B(new_n916), .C1(new_n610), .C2(new_n619), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n604), .A2(new_n607), .B1(G54), .B2(new_n527), .ZN(new_n918));
  NAND3_X1  g493(.A1(G299), .A2(new_n618), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n620), .A2(KEYINPUT105), .A3(G299), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n924), .B(KEYINPUT106), .Z(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(KEYINPUT41), .ZN(new_n926));
  OR3_X1    g501(.A1(new_n620), .A2(KEYINPUT107), .A3(G299), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n917), .A2(new_n919), .A3(KEYINPUT107), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n915), .ZN(new_n932));
  XNOR2_X1  g507(.A(G290), .B(new_n699), .ZN(new_n933));
  XNOR2_X1  g508(.A(G303), .B(new_n709), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n925), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n925), .B2(new_n932), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n849), .A2(new_n623), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(G295));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n940), .ZN(G331));
  OAI21_X1  g517(.A(G301), .B1(new_n526), .B2(new_n532), .ZN(new_n943));
  NAND4_X1  g518(.A1(G171), .A2(new_n525), .A3(new_n531), .A4(new_n529), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n857), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n857), .A3(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n945), .A2(new_n857), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n946), .A2(KEYINPUT109), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n945), .B2(new_n857), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n923), .A2(new_n951), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n931), .A2(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n935), .ZN(new_n960));
  INV_X1    g535(.A(new_n935), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n926), .A2(new_n930), .B1(new_n950), .B2(new_n952), .ZN(new_n962));
  NOR4_X1   g537(.A1(new_n954), .A2(new_n923), .A3(new_n956), .A4(new_n951), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n931), .A2(new_n953), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n957), .A2(new_n958), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n935), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n923), .A2(new_n928), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n929), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n957), .A2(new_n952), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n972), .A2(new_n973), .B1(new_n950), .B2(new_n958), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n969), .B(new_n896), .C1(new_n974), .C2(new_n935), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n966), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n964), .A2(new_n969), .A3(new_n979), .A4(new_n896), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n960), .A2(KEYINPUT110), .A3(new_n979), .A4(new_n964), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n977), .B1(new_n975), .B2(KEYINPUT43), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n978), .B1(new_n987), .B2(new_n988), .ZN(G397));
  XNOR2_X1  g564(.A(new_n803), .B(new_n806), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT112), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n786), .ZN(new_n992));
  INV_X1    g567(.A(new_n498), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n484), .B2(new_n486), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n994), .B2(new_n497), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n999), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n998), .A2(new_n1000), .B1(new_n784), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n727), .A2(new_n730), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n874), .A2(new_n731), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(G290), .B(G1986), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n997), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n1010));
  INV_X1    g585(.A(new_n996), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n499), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2078), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n499), .A2(KEYINPUT113), .A3(new_n1012), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT114), .B1(new_n995), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1023), .A2(new_n1030), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n996), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1021), .B1(new_n1032), .B2(G1961), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1022), .B(G1384), .C1(new_n994), .C2(new_n497), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n499), .B2(new_n1012), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1014), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n996), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(KEYINPUT53), .A3(new_n1018), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1010), .B1(new_n1042), .B2(G301), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT124), .B(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1017), .A2(KEYINPUT53), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1021), .B(new_n1045), .C1(new_n1032), .C2(G1961), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G171), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT126), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT50), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1031), .B1(new_n1052), .B2(new_n1027), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1011), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1054), .A2(new_n745), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(G301), .A4(new_n1045), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1055), .B2(new_n1040), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT125), .B1(new_n1046), .B2(G171), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1010), .B(new_n1057), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1981), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n582), .A2(new_n1061), .A3(new_n587), .A4(new_n592), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n513), .A2(new_n583), .ZN(new_n1063));
  AOI221_X4 g638(.A(new_n1063), .B1(new_n589), .B2(new_n591), .C1(new_n581), .C2(G651), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT117), .B(new_n1062), .C1(new_n1064), .C2(new_n1061), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n582), .A2(new_n592), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(G1981), .C1(new_n1067), .C2(new_n1063), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n1011), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1065), .A2(new_n1074), .A3(new_n1068), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n709), .A2(G1976), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(G288), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1023), .A2(new_n1011), .A3(new_n1025), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(G8), .A3(new_n1077), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1082), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT116), .B1(new_n1082), .B2(KEYINPUT52), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1076), .B(new_n1080), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G303), .A2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1011), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1072), .B2(new_n1024), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1091), .A2(G2090), .B1(G1971), .B2(new_n1017), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1092), .B2(G8), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1017), .A2(G1971), .ZN(new_n1095));
  INV_X1    g670(.A(G2090), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1011), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(KEYINPUT115), .B(new_n1097), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1101));
  OAI211_X1 g676(.A(G8), .B(new_n1088), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n996), .A2(G2084), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1966), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1107));
  OAI21_X1  g682(.A(G286), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1027), .B1(new_n1072), .B2(new_n1024), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1031), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1104), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1107), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(G168), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1108), .A2(new_n1113), .A3(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT51), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1107), .B1(new_n1053), .B2(new_n1104), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1071), .B1(new_n1116), .B2(G168), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1051), .A2(new_n1060), .A3(new_n1103), .A4(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(G299), .B(KEYINPUT57), .Z(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1089), .B1(new_n1124), .B2(KEYINPUT50), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(G1956), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1017), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1123), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1081), .A2(G2067), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1054), .B2(new_n814), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1128), .B(new_n1122), .C1(new_n1125), .C2(G1956), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n620), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(KEYINPUT122), .ZN(new_n1139));
  INV_X1    g714(.A(G1956), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1091), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n1122), .A4(new_n1128), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1139), .A2(new_n1130), .A3(new_n1143), .A4(KEYINPUT61), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1017), .A2(new_n999), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n1081), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(KEYINPUT120), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n547), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(KEYINPUT120), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n546), .B(new_n1152), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1153), .B2(new_n1150), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1138), .A2(new_n1144), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n620), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1132), .B2(KEYINPUT60), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1157), .A2(new_n1158), .B1(KEYINPUT60), .B2(new_n1132), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1135), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1121), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1085), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1093), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1116), .A2(new_n1071), .A3(G286), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1102), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1164), .A2(KEYINPUT63), .ZN(new_n1168));
  OAI21_X1  g743(.A(G8), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1088), .A2(KEYINPUT119), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI221_X1 g746(.A(G8), .B1(KEYINPUT119), .B2(new_n1088), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1168), .A2(new_n1171), .A3(new_n1162), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1094), .A2(new_n1058), .A3(new_n1102), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1118), .B1(new_n1117), .B2(new_n1108), .ZN(new_n1176));
  AOI211_X1 g751(.A(KEYINPUT51), .B(new_n1071), .C1(new_n1116), .C2(G168), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT62), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1115), .A2(new_n1179), .A3(new_n1119), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1175), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1102), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1076), .A2(new_n1078), .A3(new_n709), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1062), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1182), .A2(new_n1162), .B1(new_n1073), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1174), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1009), .B1(new_n1161), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n998), .A2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT127), .Z(new_n1190));
  OR2_X1    g765(.A1(new_n1190), .A2(KEYINPUT47), .ZN(new_n1191));
  INV_X1    g766(.A(G1986), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n735), .A2(new_n1192), .A3(new_n997), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1006), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1190), .A2(KEYINPUT47), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1002), .A2(new_n1003), .B1(G2067), .B2(new_n803), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n997), .ZN(new_n1198));
  AND4_X1   g773(.A1(new_n1191), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1187), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g775(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n696), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n906), .B2(new_n910), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n1204), .A2(new_n976), .ZN(G308));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n976), .ZN(G225));
endmodule


