

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574;

  NOR2_X2 U318 ( .A1(n420), .A2(n507), .ZN(n556) );
  XNOR2_X1 U319 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n459) );
  XNOR2_X1 U320 ( .A(KEYINPUT38), .B(n463), .ZN(n490) );
  XOR2_X1 U321 ( .A(n342), .B(n341), .Z(n286) );
  AND2_X1 U322 ( .A1(G226GAT), .A2(G233GAT), .ZN(n287) );
  NOR2_X1 U323 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U324 ( .A(n343), .B(n286), .ZN(n344) );
  XNOR2_X1 U325 ( .A(n340), .B(n287), .ZN(n313) );
  XNOR2_X1 U326 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U327 ( .A(n432), .B(n313), .ZN(n316) );
  XNOR2_X1 U328 ( .A(n460), .B(n459), .ZN(n506) );
  NOR2_X1 U329 ( .A1(n455), .A2(n437), .ZN(n552) );
  XOR2_X1 U330 ( .A(KEYINPUT41), .B(n561), .Z(n540) );
  XOR2_X1 U331 ( .A(n307), .B(n306), .Z(n520) );
  XNOR2_X1 U332 ( .A(n318), .B(n317), .ZN(n510) );
  XNOR2_X1 U333 ( .A(n438), .B(G176GAT), .ZN(n439) );
  XNOR2_X1 U334 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U335 ( .A(n440), .B(n439), .ZN(G1349GAT) );
  XNOR2_X1 U336 ( .A(n467), .B(n466), .ZN(G1328GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n289) );
  XNOR2_X1 U338 ( .A(KEYINPUT83), .B(KEYINPUT18), .ZN(n288) );
  XNOR2_X1 U339 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U340 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n291) );
  XNOR2_X1 U341 ( .A(G190GAT), .B(G183GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U343 ( .A(n293), .B(n292), .Z(n318) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n318), .B(n296), .ZN(n307) );
  XOR2_X1 U348 ( .A(G134GAT), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U349 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n297), .B(KEYINPUT81), .ZN(n406) );
  XNOR2_X1 U351 ( .A(G71GAT), .B(n406), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n301) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U356 ( .A(n303), .B(n302), .Z(n305) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G113GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  INV_X1 U359 ( .A(n520), .ZN(n455) );
  XOR2_X1 U360 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n436) );
  XOR2_X1 U361 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n309) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(G218GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U364 ( .A(G211GAT), .B(n310), .Z(n432) );
  XOR2_X1 U365 ( .A(G64GAT), .B(G204GAT), .Z(n312) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G92GAT), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n340) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(G36GAT), .ZN(n314) );
  XOR2_X1 U369 ( .A(n314), .B(G8GAT), .Z(n319) );
  INV_X1 U370 ( .A(n319), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U372 ( .A(n510), .B(KEYINPUT121), .Z(n399) );
  XNOR2_X1 U373 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n398) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G197GAT), .Z(n321) );
  XOR2_X1 U375 ( .A(G113GAT), .B(G1GAT), .Z(n410) );
  XOR2_X1 U376 ( .A(n319), .B(n410), .Z(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n326) );
  XNOR2_X1 U378 ( .A(G15GAT), .B(KEYINPUT67), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n322), .B(G22GAT), .ZN(n376) );
  XOR2_X1 U380 ( .A(n376), .B(KEYINPUT68), .Z(n324) );
  NAND2_X1 U381 ( .A1(G229GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(n326), .B(n325), .Z(n334) );
  XOR2_X1 U384 ( .A(KEYINPUT8), .B(G50GAT), .Z(n328) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G29GAT), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U387 ( .A(KEYINPUT7), .B(n329), .Z(n363) );
  XOR2_X1 U388 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n331) );
  XNOR2_X1 U389 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n363), .B(n332), .ZN(n333) );
  XOR2_X1 U392 ( .A(n334), .B(n333), .Z(n493) );
  XNOR2_X1 U393 ( .A(n493), .B(KEYINPUT69), .ZN(n548) );
  XOR2_X1 U394 ( .A(G99GAT), .B(G85GAT), .Z(n351) );
  XOR2_X1 U395 ( .A(G106GAT), .B(G78GAT), .Z(n424) );
  XNOR2_X1 U396 ( .A(n351), .B(n424), .ZN(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n336) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n380) );
  XOR2_X1 U400 ( .A(KEYINPUT33), .B(n380), .Z(n338) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n345) );
  XNOR2_X1 U403 ( .A(G120GAT), .B(G57GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n339), .B(G148GAT), .ZN(n405) );
  XNOR2_X1 U405 ( .A(n340), .B(n405), .ZN(n343) );
  XOR2_X1 U406 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n342) );
  XNOR2_X1 U407 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n341) );
  XOR2_X1 U408 ( .A(n347), .B(n346), .Z(n561) );
  INV_X1 U409 ( .A(n561), .ZN(n461) );
  XOR2_X1 U410 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n386) );
  XOR2_X1 U411 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n349) );
  NAND2_X1 U412 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U414 ( .A(KEYINPUT74), .B(n350), .ZN(n361) );
  XOR2_X1 U415 ( .A(G106GAT), .B(G162GAT), .Z(n353) );
  XOR2_X1 U416 ( .A(G134GAT), .B(KEYINPUT76), .Z(n409) );
  XNOR2_X1 U417 ( .A(n351), .B(n409), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U419 ( .A(n354), .B(G218GAT), .Z(n359) );
  XOR2_X1 U420 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n356) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U423 ( .A(G190GAT), .B(n357), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n468) );
  XNOR2_X1 U427 ( .A(n468), .B(KEYINPUT99), .ZN(n364) );
  XNOR2_X1 U428 ( .A(KEYINPUT36), .B(n364), .ZN(n569) );
  XOR2_X1 U429 ( .A(G211GAT), .B(KEYINPUT79), .Z(n366) );
  XNOR2_X1 U430 ( .A(G183GAT), .B(KEYINPUT77), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n384) );
  XOR2_X1 U432 ( .A(KEYINPUT80), .B(G57GAT), .Z(n368) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(G1GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n370) );
  XNOR2_X1 U436 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U438 ( .A(n372), .B(n371), .Z(n378) );
  XOR2_X1 U439 ( .A(G64GAT), .B(G78GAT), .Z(n374) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U444 ( .A(n379), .B(G155GAT), .Z(n382) );
  XNOR2_X1 U445 ( .A(G127GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n565) );
  NAND2_X1 U448 ( .A1(n569), .A2(n565), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n387) );
  NAND2_X1 U450 ( .A1(n461), .A2(n387), .ZN(n388) );
  NOR2_X1 U451 ( .A1(n548), .A2(n388), .ZN(n389) );
  XNOR2_X1 U452 ( .A(KEYINPUT111), .B(n389), .ZN(n396) );
  XOR2_X1 U453 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n391) );
  INV_X1 U454 ( .A(n493), .ZN(n557) );
  NAND2_X1 U455 ( .A1(n557), .A2(n540), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n393) );
  INV_X1 U457 ( .A(n565), .ZN(n469) );
  NAND2_X1 U458 ( .A1(n469), .A2(n468), .ZN(n392) );
  XNOR2_X1 U459 ( .A(KEYINPUT47), .B(n394), .ZN(n395) );
  NAND2_X1 U460 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n517) );
  NAND2_X1 U462 ( .A1(n399), .A2(n517), .ZN(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT54), .B(n400), .ZN(n420) );
  XNOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n401), .B(KEYINPUT88), .ZN(n402) );
  XOR2_X1 U466 ( .A(n402), .B(KEYINPUT2), .Z(n404) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(G162GAT), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n431) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n418) );
  XOR2_X1 U470 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n408) );
  XNOR2_X1 U471 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n414) );
  XOR2_X1 U473 ( .A(n409), .B(G85GAT), .Z(n412) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U476 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n431), .B(n419), .ZN(n448) );
  XNOR2_X1 U481 ( .A(KEYINPUT89), .B(n448), .ZN(n507) );
  XOR2_X1 U482 ( .A(G148GAT), .B(G204GAT), .Z(n422) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(G22GAT), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U485 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U488 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n428) );
  XNOR2_X1 U489 ( .A(KEYINPUT22), .B(KEYINPUT86), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U491 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n450) );
  NAND2_X1 U494 ( .A1(n556), .A2(n450), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U496 ( .A1(n552), .A2(n540), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT90), .B(KEYINPUT27), .Z(n441) );
  XOR2_X1 U499 ( .A(n510), .B(n441), .Z(n451) );
  NOR2_X1 U500 ( .A1(n520), .A2(n450), .ZN(n442) );
  XOR2_X1 U501 ( .A(n442), .B(KEYINPUT26), .Z(n537) );
  INV_X1 U502 ( .A(n537), .ZN(n555) );
  NAND2_X1 U503 ( .A1(n451), .A2(n555), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n443), .B(KEYINPUT92), .ZN(n447) );
  NAND2_X1 U505 ( .A1(n510), .A2(n520), .ZN(n444) );
  NAND2_X1 U506 ( .A1(n450), .A2(n444), .ZN(n445) );
  XOR2_X1 U507 ( .A(KEYINPUT25), .B(n445), .Z(n446) );
  NAND2_X1 U508 ( .A1(n447), .A2(n446), .ZN(n449) );
  NAND2_X1 U509 ( .A1(n449), .A2(n448), .ZN(n457) );
  XOR2_X1 U510 ( .A(n450), .B(KEYINPUT28), .Z(n519) );
  NAND2_X1 U511 ( .A1(n451), .A2(n507), .ZN(n452) );
  XNOR2_X1 U512 ( .A(KEYINPUT91), .B(n452), .ZN(n518) );
  INV_X1 U513 ( .A(n518), .ZN(n453) );
  NOR2_X1 U514 ( .A1(n519), .A2(n453), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n457), .A2(n456), .ZN(n471) );
  NAND2_X1 U517 ( .A1(n569), .A2(n471), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n458), .A2(n565), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n548), .A2(n461), .ZN(n473) );
  NOR2_X1 U520 ( .A1(n506), .A2(n473), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT101), .B(n462), .Z(n463) );
  NAND2_X1 U522 ( .A1(n507), .A2(n490), .ZN(n467) );
  XOR2_X1 U523 ( .A(G29GAT), .B(KEYINPUT102), .Z(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT34), .B(KEYINPUT93), .Z(n475) );
  INV_X1 U526 ( .A(n468), .ZN(n551) );
  NOR2_X1 U527 ( .A1(n551), .A2(n469), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT16), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n494) );
  NOR2_X1 U530 ( .A1(n473), .A2(n494), .ZN(n484) );
  NAND2_X1 U531 ( .A1(n484), .A2(n507), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n478) );
  NAND2_X1 U535 ( .A1(n484), .A2(n510), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT35), .B(KEYINPUT97), .Z(n481) );
  NAND2_X1 U539 ( .A1(n484), .A2(n520), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n483) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT96), .Z(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n484), .A2(n519), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(KEYINPUT98), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  NAND2_X1 U546 ( .A1(n490), .A2(n510), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U548 ( .A1(n490), .A2(n520), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NAND2_X1 U551 ( .A1(n490), .A2(n519), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G50GAT), .B(n492), .ZN(G1331GAT) );
  NAND2_X1 U554 ( .A1(n493), .A2(n540), .ZN(n505) );
  NOR2_X1 U555 ( .A1(n505), .A2(n494), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT105), .B(n495), .Z(n502) );
  NAND2_X1 U557 ( .A1(n502), .A2(n507), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1332GAT) );
  NAND2_X1 U561 ( .A1(n502), .A2(n510), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U563 ( .A(G71GAT), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U564 ( .A1(n502), .A2(n520), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(G78GAT), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U567 ( .A1(n502), .A2(n519), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  XNOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n509) );
  NOR2_X1 U570 ( .A1(n506), .A2(n505), .ZN(n513) );
  NAND2_X1 U571 ( .A1(n507), .A2(n513), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NAND2_X1 U573 ( .A1(n513), .A2(n510), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U575 ( .A1(n520), .A2(n513), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n515) );
  NAND2_X1 U578 ( .A1(n513), .A2(n519), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  XNOR2_X1 U581 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n536) );
  NOR2_X1 U583 ( .A1(n519), .A2(n536), .ZN(n521) );
  NAND2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT113), .B(n522), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n548), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT49), .Z(n526) );
  NAND2_X1 U589 ( .A1(n532), .A2(n540), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n528) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(n529), .Z(n531) );
  NAND2_X1 U595 ( .A1(n532), .A2(n565), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U598 ( .A1(n532), .A2(n551), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U602 ( .A(KEYINPUT119), .B(n538), .Z(n545) );
  NAND2_X1 U603 ( .A1(n545), .A2(n557), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  NAND2_X1 U606 ( .A1(n545), .A2(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n565), .A2(n545), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n551), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G162GAT), .B(n547), .ZN(G1347GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n552), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G169GAT), .B(n549), .ZN(G1348GAT) );
  NAND2_X1 U616 ( .A1(n565), .A2(n552), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT58), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G190GAT), .B(n554), .ZN(G1351GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n559) );
  AND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n570), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G197GAT), .B(n560), .ZN(G1352GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n563) );
  NAND2_X1 U627 ( .A1(n570), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G204GAT), .B(n564), .Z(G1353GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n567) );
  NAND2_X1 U631 ( .A1(n570), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G211GAT), .B(n568), .ZN(G1354GAT) );
  XNOR2_X1 U634 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1355GAT) );
endmodule

