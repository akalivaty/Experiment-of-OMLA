//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT25), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n187), .A2(KEYINPUT25), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n196), .B2(new_n190), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n200), .A2(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n203), .C1(new_n204), .C2(KEYINPUT23), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT24), .B(G110), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(G119), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(new_n201), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n205), .A2(G110), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(new_n210), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n197), .A2(new_n198), .ZN(new_n212));
  XNOR2_X1  g026(.A(G125), .B(G140), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n214), .B2(new_n213), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n205), .A2(G110), .B1(new_n207), .B2(new_n209), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT22), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(G137), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n219), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G902), .ZN(new_n225));
  AOI211_X1 g039(.A(new_n188), .B(new_n189), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n188), .ZN(new_n227));
  INV_X1    g041(.A(G234), .ZN(new_n228));
  OAI21_X1  g042(.A(G217), .B1(new_n228), .B2(G902), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT73), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n225), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n224), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT20), .ZN(new_n237));
  INV_X1    g051(.A(G131), .ZN(new_n238));
  INV_X1    g052(.A(G237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n220), .A3(G214), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n239), .A2(new_n220), .A3(G143), .A4(G214), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT17), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n197), .B(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n243), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n245), .B(new_n246), .C1(new_n249), .C2(KEYINPUT17), .ZN(new_n250));
  XNOR2_X1  g064(.A(G113), .B(G122), .ZN(new_n251));
  INV_X1    g065(.A(G104), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n242), .A2(new_n254), .A3(new_n243), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT18), .A2(G131), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n216), .B1(new_n198), .B2(new_n213), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT87), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT87), .B1(new_n257), .B2(new_n258), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n250), .B(new_n253), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n212), .B1(new_n244), .B2(new_n248), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT88), .B1(new_n213), .B2(new_n214), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT19), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n265), .B2(new_n264), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n263), .A2(new_n264), .B1(new_n213), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n257), .A2(new_n258), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT87), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT87), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n261), .B1(new_n274), .B2(new_n253), .ZN(new_n275));
  NOR2_X1   g089(.A1(G475), .A2(G902), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n237), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n237), .A3(new_n276), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n273), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n253), .B1(new_n281), .B2(new_n250), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n282), .B2(KEYINPUT89), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n250), .B1(new_n259), .B2(new_n260), .ZN(new_n284));
  INV_X1    g098(.A(new_n253), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT89), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n261), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G475), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n280), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G128), .B(G143), .ZN(new_n292));
  INV_X1    g106(.A(G134), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT77), .B(G107), .ZN(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G122), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G107), .ZN(new_n298));
  INV_X1    g112(.A(G122), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n300), .B2(KEYINPUT14), .ZN(new_n301));
  XOR2_X1   g115(.A(G116), .B(G122), .Z(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(KEYINPUT14), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n294), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n295), .B(new_n296), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n292), .A2(KEYINPUT13), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n202), .A2(KEYINPUT13), .A3(G143), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n293), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n306), .A2(new_n308), .B1(new_n293), .B2(new_n292), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n312), .A2(new_n313), .A3(G953), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT91), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n304), .A2(new_n310), .A3(new_n314), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n317), .B(new_n319), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G478), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n325), .A2(KEYINPUT15), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n324), .A2(new_n225), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n324), .B2(new_n225), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n291), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G952), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G953), .ZN(new_n333));
  NAND2_X1  g147(.A1(G234), .A2(G237), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n335), .B(KEYINPUT92), .Z(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(G902), .A3(G953), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT21), .B(G898), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n343));
  NOR2_X1   g157(.A1(G472), .A2(G902), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n293), .A2(G137), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(KEYINPUT11), .ZN(new_n348));
  INV_X1    g162(.A(G137), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT11), .B1(new_n349), .B2(G134), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT67), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(KEYINPUT11), .A3(G134), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(KEYINPUT68), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n349), .A2(G134), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n355), .B2(KEYINPUT68), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G131), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n351), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(new_n238), .A3(new_n354), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n241), .A2(G146), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT65), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n241), .A2(KEYINPUT65), .A3(G146), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n198), .A2(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT0), .A2(G128), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR3_X1   g184(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n367), .A2(new_n362), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n368), .A2(new_n374), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n361), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n378), .A3(G128), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n364), .A2(new_n365), .B1(G143), .B2(new_n198), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n202), .B1(new_n367), .B2(KEYINPUT1), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G131), .B1(new_n347), .B2(new_n355), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n360), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(KEYINPUT30), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n386));
  INV_X1    g200(.A(G116), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(G119), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n200), .A2(KEYINPUT69), .A3(G116), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n388), .A2(new_n389), .B1(new_n387), .B2(G119), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT2), .B(G113), .Z(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT70), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n382), .A2(new_n360), .A3(new_n383), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT66), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n375), .A2(new_n370), .ZN(new_n402));
  INV_X1    g216(.A(new_n373), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n369), .B1(new_n403), .B2(new_n371), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n380), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n358), .A2(new_n360), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n376), .A2(KEYINPUT66), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n385), .B(new_n399), .C1(new_n408), .C2(KEYINPUT30), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n400), .B1(new_n361), .B2(new_n376), .ZN(new_n410));
  INV_X1    g224(.A(new_n399), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n239), .A2(new_n220), .A3(G210), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT26), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(G101), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT71), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n409), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT31), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n409), .A2(new_n418), .A3(KEYINPUT31), .A4(new_n412), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n410), .A2(KEYINPUT28), .A3(new_n411), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(new_n426), .C1(new_n411), .C2(new_n408), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n345), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n343), .B1(new_n429), .B2(KEYINPUT72), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT72), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n421), .A2(new_n422), .B1(new_n427), .B2(new_n417), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n431), .B(KEYINPUT32), .C1(new_n432), .C2(new_n345), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n410), .A2(new_n411), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n425), .A2(new_n426), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n417), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT29), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n412), .A2(new_n417), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n427), .A2(new_n437), .B1(new_n409), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n225), .B(new_n438), .C1(new_n440), .C2(KEYINPUT29), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G472), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n236), .B(new_n342), .C1(new_n434), .C2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G214), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n379), .B(new_n194), .C1(new_n380), .C2(new_n381), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(KEYINPUT85), .C1(new_n376), .C2(new_n194), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n405), .A2(new_n448), .A3(G125), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G224), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G953), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n447), .B(new_n449), .C1(new_n451), .C2(G953), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n452), .A2(KEYINPUT7), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n450), .A2(KEYINPUT7), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G122), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n459), .B(KEYINPUT8), .Z(new_n460));
  NAND2_X1  g274(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n200), .A2(G116), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(G113), .C1(KEYINPUT5), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n392), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n298), .A2(KEYINPUT77), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT77), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G107), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n467), .A3(G104), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT78), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT76), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT76), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT78), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n295), .A3(new_n476), .A4(G104), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(new_n252), .B2(G107), .ZN(new_n478));
  AOI21_X1  g292(.A(G101), .B1(new_n252), .B2(G107), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n470), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n295), .A2(G104), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n252), .A2(G107), .ZN(new_n482));
  OAI21_X1  g296(.A(G101), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n483), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n464), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n464), .A2(new_n484), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n460), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n458), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n252), .A2(G107), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n470), .A2(new_n477), .A3(new_n493), .A4(new_n478), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n494), .A2(G101), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n480), .A2(KEYINPUT4), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(KEYINPUT79), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT79), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n480), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(G101), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(new_n503), .A3(G101), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n399), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n489), .B(new_n459), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n492), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n459), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n499), .A2(new_n498), .A3(new_n500), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT79), .B1(new_n495), .B2(new_n496), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n512), .B2(new_n488), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n506), .A3(KEYINPUT6), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n453), .A2(new_n454), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(new_n509), .C1(new_n512), .C2(new_n488), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G210), .B1(G237), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n507), .A2(new_n518), .A3(new_n520), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n445), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n525));
  INV_X1    g339(.A(G469), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G140), .ZN(new_n527));
  INV_X1    g341(.A(G227), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(G953), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n527), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n361), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n483), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT80), .B1(new_n480), .B2(new_n483), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(new_n536), .A3(new_n382), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n480), .A2(new_n483), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n379), .B1(new_n375), .B2(new_n381), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n534), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n382), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n486), .A2(new_n547), .A3(new_n487), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n539), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n544), .A3(new_n534), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n553));
  AND4_X1   g367(.A1(new_n553), .A2(new_n480), .A3(new_n539), .A4(new_n483), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n547), .B1(new_n486), .B2(new_n487), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(new_n553), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n504), .A2(new_n376), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n497), .B2(new_n501), .ZN(new_n560));
  INV_X1    g374(.A(new_n361), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n531), .B1(new_n552), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n382), .B1(new_n535), .B2(new_n536), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n554), .B1(new_n564), .B2(KEYINPUT10), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n558), .B1(new_n511), .B2(new_n510), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n361), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n567), .A2(new_n562), .A3(new_n531), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT82), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n544), .B1(new_n550), .B2(new_n534), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n545), .B(new_n533), .C1(new_n548), .C2(new_n549), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n565), .A2(new_n566), .A3(new_n361), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n530), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n567), .A2(new_n562), .A3(new_n531), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n526), .B1(new_n578), .B2(new_n225), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n567), .A2(new_n562), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n530), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n552), .A2(new_n562), .A3(new_n531), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT83), .B(G469), .Z(new_n584));
  AND3_X1   g398(.A1(new_n583), .A2(new_n225), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n524), .B(new_n525), .C1(new_n579), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n443), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(new_n429), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n432), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n236), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n525), .C1(new_n579), .C2(new_n585), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n275), .A2(new_n237), .A3(new_n276), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n277), .ZN(new_n597));
  INV_X1    g411(.A(G475), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n283), .B2(new_n288), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n314), .A2(KEYINPUT95), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n311), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT33), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n324), .B2(KEYINPUT33), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n325), .A2(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n324), .A2(new_n225), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT96), .B(G478), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n522), .A2(KEYINPUT94), .A3(new_n523), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n507), .A2(new_n518), .A3(new_n612), .A4(new_n520), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n613), .A2(new_n444), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NOR4_X1   g429(.A1(new_n595), .A2(new_n340), .A3(new_n610), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n595), .ZN(new_n619));
  NOR4_X1   g433(.A1(new_n597), .A2(new_n599), .A3(new_n329), .A4(new_n340), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n611), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT35), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G107), .ZN(G9));
  INV_X1    g439(.A(new_n223), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n219), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n234), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n226), .B2(new_n231), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n342), .A2(new_n593), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n587), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  NAND2_X1  g449(.A1(new_n613), .A2(new_n444), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n507), .A2(new_n518), .A3(new_n520), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n520), .B1(new_n507), .B2(new_n518), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n639), .B2(KEYINPUT94), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n434), .A2(new_n442), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n600), .A2(new_n330), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n337), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n336), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n525), .B(new_n630), .C1(new_n579), .C2(new_n585), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n202), .ZN(G30));
  NOR4_X1   g464(.A1(new_n600), .A2(new_n630), .A3(new_n445), .A4(new_n329), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n639), .B(KEYINPUT38), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n439), .B2(new_n435), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n409), .A2(new_n412), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n437), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n430), .A2(new_n433), .B1(G472), .B2(new_n657), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n652), .A2(new_n653), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n525), .B1(new_n579), .B2(new_n585), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n645), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n661), .A2(KEYINPUT40), .A3(new_n662), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n659), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n241), .ZN(G45));
  NOR3_X1   g482(.A1(new_n600), .A2(new_n608), .A3(new_n645), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n640), .A2(new_n641), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n648), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n198), .ZN(G48));
  AOI21_X1  g486(.A(new_n236), .B1(new_n434), .B2(new_n442), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n340), .B(new_n608), .C1(new_n280), .C2(new_n290), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n583), .A2(new_n225), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n583), .A2(new_n225), .A3(new_n584), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n525), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n640), .A3(new_n674), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  NAND3_X1  g496(.A1(new_n621), .A2(new_n673), .A3(new_n679), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  INV_X1    g498(.A(new_n342), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n641), .A2(new_n685), .A3(new_n630), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n640), .A2(new_n679), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT99), .B1(new_n615), .B2(new_n678), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n200), .ZN(G21));
  OAI21_X1  g506(.A(new_n423), .B1(new_n437), .B2(new_n436), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n344), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n592), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n340), .A3(new_n236), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n600), .A2(new_n329), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n640), .A3(new_n679), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT101), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  NOR2_X1   g514(.A1(new_n695), .A2(new_n631), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n669), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n688), .B2(new_n689), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n194), .ZN(G27));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n574), .A2(new_n576), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n526), .B1(new_n706), .B2(new_n225), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n705), .B1(new_n585), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n574), .B2(new_n576), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n677), .B(KEYINPUT102), .C1(new_n526), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n522), .A2(new_n523), .ZN(new_n712));
  INV_X1    g526(.A(new_n525), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n445), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OR3_X1    g529(.A1(new_n429), .A2(KEYINPUT104), .A3(KEYINPUT32), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n429), .B2(KEYINPUT32), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n716), .A2(new_n442), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n669), .A2(KEYINPUT42), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n235), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n673), .A2(new_n711), .A3(new_n714), .A4(new_n669), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n723));
  AOI22_X1  g537(.A1(new_n715), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n238), .ZN(G33));
  NAND4_X1  g539(.A1(new_n673), .A2(new_n711), .A3(new_n714), .A4(new_n646), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n526), .A2(new_n225), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n706), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n526), .B1(new_n578), .B2(new_n731), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(KEYINPUT105), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n569), .B2(new_n577), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n735), .B1(new_n736), .B2(new_n526), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT106), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n563), .A2(new_n568), .A3(KEYINPUT82), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n731), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .A3(G469), .ZN(new_n742));
  INV_X1    g556(.A(new_n732), .ZN(new_n743));
  AND4_X1   g557(.A1(KEYINPUT106), .A2(new_n742), .A3(new_n737), .A4(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n730), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n737), .A3(new_n743), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n734), .A2(KEYINPUT106), .A3(new_n737), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n730), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n585), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n662), .A2(new_n525), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n728), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n752), .B1(new_n751), .B2(new_n730), .ZN(new_n757));
  AOI211_X1 g571(.A(KEYINPUT46), .B(new_n729), .C1(new_n749), .C2(new_n750), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n677), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n755), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(KEYINPUT107), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n608), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n600), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT43), .Z(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n593), .A3(new_n630), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n712), .A2(new_n445), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n756), .A2(new_n761), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT108), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  OAI21_X1  g588(.A(KEYINPUT47), .B1(new_n754), .B2(new_n713), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n759), .A2(new_n776), .A3(new_n525), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n669), .A2(new_n236), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n770), .A2(new_n641), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  INV_X1    g595(.A(new_n336), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n764), .A2(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n236), .A3(new_n695), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n445), .A3(new_n653), .A4(new_n679), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT50), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n783), .A2(new_n678), .A3(new_n770), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n701), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n236), .A2(new_n336), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n679), .A2(new_n769), .A3(new_n658), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n600), .A2(new_n608), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT116), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(KEYINPUT116), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n676), .A2(new_n677), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n525), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n775), .B2(new_n777), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n784), .A2(new_n769), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n797), .B(KEYINPUT115), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n754), .A2(KEYINPUT47), .A3(new_n713), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n776), .B1(new_n759), .B2(new_n525), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n799), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n792), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n800), .A2(KEYINPUT51), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n648), .B1(new_n647), .B2(new_n670), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n703), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n658), .A2(new_n713), .A3(new_n630), .A4(new_n645), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n615), .A2(new_n329), .A3(new_n600), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n711), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n688), .A2(new_n689), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n592), .A2(new_n669), .A3(new_n630), .A4(new_n694), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n615), .B1(new_n434), .B2(new_n442), .ZN(new_n818));
  INV_X1    g632(.A(new_n648), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n818), .B(new_n819), .C1(new_n646), .C2(new_n669), .ZN(new_n820));
  AND4_X1   g634(.A1(KEYINPUT52), .A2(new_n817), .A3(new_n820), .A4(new_n813), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n680), .A2(new_n683), .A3(new_n698), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n724), .A2(new_n690), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n711), .A3(new_n714), .ZN(new_n825));
  INV_X1    g639(.A(new_n645), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n641), .A2(new_n769), .A3(new_n331), .A4(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n726), .B(new_n825), .C1(new_n648), .C2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n620), .B(new_n444), .C1(new_n637), .C2(new_n638), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n712), .A2(new_n444), .A3(new_n674), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT110), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n524), .A2(new_n834), .A3(new_n674), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n595), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n673), .A2(new_n341), .A3(new_n331), .ZN(new_n838));
  INV_X1    g652(.A(new_n632), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n586), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n828), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n824), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n822), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n823), .A2(new_n690), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n721), .A2(new_n715), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n722), .A2(new_n723), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n726), .A2(new_n825), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n827), .A2(new_n648), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n833), .A2(new_n835), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n829), .B(KEYINPUT111), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n619), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n587), .B1(new_n443), .B2(new_n632), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n844), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n824), .A2(new_n841), .A3(KEYINPUT112), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n817), .A2(new_n820), .A3(new_n813), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n810), .A2(KEYINPUT52), .A3(new_n813), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT113), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n814), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n843), .B(KEYINPUT54), .C1(new_n861), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n724), .A2(new_n823), .A3(new_n871), .A4(new_n690), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n855), .A4(new_n856), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n849), .A2(new_n871), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n868), .A3(new_n866), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n859), .B1(new_n822), .B2(new_n842), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n719), .A2(new_n235), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n787), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n882));
  OR2_X1    g696(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI221_X1 g698(.A(new_n333), .B1(new_n790), .B2(new_n610), .C1(new_n881), .C2(new_n882), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n884), .B(new_n885), .C1(new_n815), .C2(new_n784), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n870), .A2(new_n879), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT118), .B1(new_n808), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n870), .A2(new_n879), .A3(new_n886), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n802), .A2(new_n803), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n805), .B1(new_n892), .B2(new_n797), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(new_n795), .ZN(new_n894));
  INV_X1    g708(.A(new_n807), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n804), .B2(new_n805), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n889), .B(new_n890), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n332), .A2(new_n220), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n888), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n236), .A2(new_n763), .A3(new_n713), .A4(new_n445), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT109), .Z(new_n901));
  XOR2_X1   g715(.A(new_n796), .B(KEYINPUT49), .Z(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n653), .A3(new_n658), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(G75));
  NOR2_X1   g718(.A1(new_n220), .A2(G952), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n873), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n845), .A2(KEYINPUT114), .A3(new_n848), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n875), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n869), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n842), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n864), .A2(new_n865), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT53), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n225), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n514), .A2(new_n517), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n515), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n906), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n915), .A2(G210), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G51));
  AOI211_X1 g740(.A(new_n225), .B(new_n751), .C1(new_n876), .C2(new_n878), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n729), .B(KEYINPUT57), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n927), .B1(new_n931), .B2(new_n583), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT120), .B1(new_n932), .B2(new_n905), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT120), .ZN(new_n934));
  INV_X1    g748(.A(new_n583), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT54), .B1(new_n910), .B2(new_n913), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n879), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n934), .B(new_n906), .C1(new_n938), .C2(new_n927), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n933), .A2(new_n939), .ZN(G54));
  NAND3_X1  g754(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  INV_X1    g755(.A(new_n275), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n905), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .A4(new_n275), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(G60));
  XNOR2_X1  g759(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n325), .A2(new_n225), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n870), .B2(new_n879), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n906), .B1(new_n950), .B2(new_n604), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n604), .A2(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n936), .B2(new_n879), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(G63));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n914), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n628), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n224), .B(KEYINPUT123), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n906), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n957), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n960), .A2(new_n963), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n961), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(G66));
  NAND2_X1  g782(.A1(new_n855), .A2(new_n856), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n969), .A2(new_n690), .A3(new_n823), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n220), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n338), .B2(new_n451), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n917), .B1(G898), .B2(new_n220), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  AOI21_X1  g791(.A(new_n220), .B1(G227), .B2(G900), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n610), .A2(new_n642), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n673), .A2(new_n769), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n663), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n810), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n667), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n667), .B2(new_n983), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n772), .A3(new_n780), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n385), .B1(new_n408), .B2(KEYINPUT30), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(new_n267), .Z(new_n990));
  AND3_X1   g804(.A1(new_n988), .A2(new_n220), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n880), .A2(new_n812), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n756), .A2(new_n761), .A3(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n810), .A2(new_n848), .A3(new_n726), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n772), .A2(new_n780), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n995), .B2(new_n220), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n979), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n990), .A2(new_n528), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n998), .B2(new_n643), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(new_n439), .A2(new_n409), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  AND3_X1   g817(.A1(new_n656), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n843), .B(new_n1004), .C1(new_n861), .C2(new_n869), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n987), .A2(new_n772), .A3(new_n780), .A4(new_n970), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1007), .A2(new_n1003), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n1008), .B2(new_n656), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n780), .A2(new_n993), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n772), .A2(new_n994), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n970), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1001), .B1(new_n1013), .B2(new_n1003), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1014), .B2(new_n905), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1003), .B1(new_n995), .B2(new_n971), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n409), .A3(new_n439), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1017), .A2(KEYINPUT126), .A3(new_n906), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1009), .B1(new_n1015), .B2(new_n1018), .ZN(G57));
endmodule


