//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G228gat), .A2(G233gat), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n208), .B(KEYINPUT78), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT29), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G211gat), .A2(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT22), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT71), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT71), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n212), .B2(new_n213), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n219), .B(new_n211), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n210), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT73), .B(KEYINPUT3), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT2), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237));
  NAND2_X1  g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n246));
  INV_X1    g045(.A(new_n211), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n223), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n243), .A3(new_n226), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n210), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n209), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n235), .A2(new_n243), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT3), .B1(new_n225), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT29), .B1(new_n248), .B2(new_n223), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT79), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n251), .A2(new_n210), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n249), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n250), .A2(KEYINPUT80), .A3(new_n252), .ZN(new_n264));
  INV_X1    g063(.A(new_n208), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n254), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT81), .B1(new_n260), .B2(new_n266), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n207), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT3), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n258), .B2(KEYINPUT79), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n225), .A2(new_n256), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n244), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n208), .B1(new_n253), .B2(new_n261), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n275), .A2(new_n268), .A3(new_n264), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n254), .ZN(new_n278));
  AND4_X1   g077(.A1(new_n270), .A2(new_n277), .A3(new_n278), .A4(new_n207), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n204), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n269), .A2(KEYINPUT82), .A3(new_n206), .A4(new_n270), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n270), .A2(new_n277), .A3(new_n206), .A4(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n277), .A3(new_n278), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G22gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n204), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT84), .B(new_n204), .C1(new_n271), .C2(new_n279), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G227gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT64), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(G169gat), .A3(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT23), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(KEYINPUT23), .ZN(new_n312));
  AND4_X1   g111(.A1(new_n304), .A2(new_n309), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(KEYINPUT23), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT65), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n315), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n312), .ZN(new_n322));
  OAI22_X1  g121(.A1(new_n313), .A2(KEYINPUT25), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n306), .A2(new_n308), .B1(new_n326), .B2(KEYINPUT26), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n317), .A2(new_n328), .A3(new_n318), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT68), .A3(new_n301), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT27), .B(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT28), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n336), .A2(new_n338), .A3(new_n333), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n339), .B2(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT68), .B1(new_n330), .B2(new_n301), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n323), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G113gat), .B(G120gat), .ZN(new_n344));
  INV_X1    g143(.A(G127gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(G134gat), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G127gat), .ZN(new_n348));
  OAI22_X1  g147(.A1(new_n344), .A2(KEYINPUT1), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G120gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G113gat), .ZN(new_n351));
  INV_X1    g150(.A(G113gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G120gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G127gat), .B(G134gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT69), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n343), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n359), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n330), .A2(new_n301), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n331), .A3(new_n340), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n368), .B2(new_n323), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n299), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n296), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n299), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n343), .A2(new_n362), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n364), .A3(new_n323), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT70), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n370), .A2(new_n379), .A3(KEYINPUT32), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n374), .A2(new_n373), .A3(new_n375), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n382), .B(KEYINPUT34), .Z(new_n383));
  OAI211_X1 g182(.A(new_n370), .B(KEYINPUT32), .C1(new_n371), .C2(new_n296), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n381), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT87), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n293), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n343), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n368), .A2(G226gat), .A3(G233gat), .A4(new_n323), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n249), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n397), .A3(new_n249), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n402), .ZN(new_n405));
  INV_X1    g204(.A(new_n403), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT30), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(new_n405), .C1(new_n406), .C2(new_n398), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT72), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n251), .A2(new_n358), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n244), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n359), .A2(new_n429), .A3(new_n255), .A4(new_n361), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n349), .A2(new_n357), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n255), .A3(KEYINPUT74), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n358), .B2(new_n244), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT76), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n430), .A2(new_n436), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n423), .B(new_n428), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n432), .A2(new_n434), .B1(new_n244), .B2(new_n358), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n419), .B1(new_n440), .B2(new_n420), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n429), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n427), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n362), .A2(new_n244), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n421), .B1(new_n446), .B2(KEYINPUT4), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n417), .B1(new_n439), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n428), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n422), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n444), .A3(new_n443), .ZN(new_n452));
  INV_X1    g251(.A(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n416), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n449), .A2(new_n455), .A3(KEYINPUT86), .A4(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n449), .B2(new_n456), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n416), .B1(new_n451), .B2(new_n454), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT77), .A3(KEYINPUT6), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(KEYINPUT6), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT86), .B1(new_n463), .B2(new_n455), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n411), .B(new_n412), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT89), .B1(new_n394), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n387), .A2(new_n393), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n411), .A2(new_n412), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n455), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n468), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n467), .A2(new_n473), .A3(new_n474), .A4(new_n293), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n385), .A2(new_n386), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n293), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n411), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n459), .A2(new_n461), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n470), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n481), .A2(new_n293), .ZN(new_n485));
  OR3_X1    g284(.A1(new_n450), .A2(KEYINPUT39), .A3(new_n420), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n440), .B2(new_n420), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n450), .B2(new_n420), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT40), .A4(new_n416), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT85), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n489), .A2(new_n416), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT40), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n493), .A2(new_n411), .A3(new_n460), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n399), .A2(new_n496), .A3(new_n403), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT37), .B1(new_n406), .B2(new_n398), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT38), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n499), .A2(new_n402), .B1(new_n500), .B2(new_n407), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT38), .B(new_n405), .C1(new_n497), .C2(new_n498), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n469), .A2(new_n472), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n495), .A2(new_n504), .A3(new_n293), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n477), .B(KEYINPUT36), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n484), .B1(new_n485), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(G169gat), .B(G197gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT12), .Z(new_n514));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(G1gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  MUX2_X1   g317(.A(G1gat), .B(new_n517), .S(new_n518), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G8gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT91), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT92), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT92), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT14), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n522), .A2(KEYINPUT15), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n522), .A2(KEYINPUT94), .A3(KEYINPUT15), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n521), .A2(KEYINPUT15), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n520), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n533), .A2(new_n540), .A3(new_n520), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n515), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(KEYINPUT96), .B(new_n547), .C1(new_n542), .C2(new_n543), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n533), .A2(new_n540), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n533), .B2(new_n540), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n520), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n546), .A3(new_n542), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n549), .A2(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n540), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT17), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n533), .A2(new_n540), .A3(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n541), .B1(new_n561), .B2(new_n520), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT18), .B1(new_n562), .B2(new_n546), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n514), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n548), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT96), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n515), .A3(new_n548), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(KEYINPUT18), .A3(new_n546), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n555), .A2(new_n556), .ZN(new_n570));
  INV_X1    g369(.A(new_n514), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n564), .A2(KEYINPUT97), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT97), .B1(new_n564), .B2(new_n572), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n508), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n520), .ZN(new_n578));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n578), .B1(KEYINPUT21), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT98), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(new_n595), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n587), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n593), .A2(new_n595), .ZN(new_n599));
  INV_X1    g398(.A(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G183gat), .B(G211gat), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n598), .B2(new_n602), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT99), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT100), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(KEYINPUT8), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT101), .B(G85gat), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n617), .B(new_n618), .C1(G92gat), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n559), .B2(new_n560), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n558), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n614), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n622), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n552), .B2(new_n553), .ZN(new_n629));
  INV_X1    g428(.A(new_n614), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n629), .A2(new_n625), .A3(new_n624), .A4(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n613), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n631), .A3(new_n611), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT103), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT104), .B1(new_n607), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n598), .A2(new_n602), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n603), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n635), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n631), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n633), .B1(new_n645), .B2(new_n612), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT102), .B(new_n613), .C1(new_n627), .C2(new_n631), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n638), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n622), .B(new_n585), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT105), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n586), .A2(new_n622), .A3(new_n658), .A4(KEYINPUT10), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G120gat), .B(G148gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT106), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n663), .B(new_n668), .C1(new_n653), .C2(new_n662), .ZN(new_n669));
  INV_X1    g468(.A(new_n662), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n655), .B2(new_n660), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n653), .A2(new_n662), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n652), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n577), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n470), .A2(new_n461), .A3(new_n459), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(G1gat), .Z(G1324gat));
  OAI21_X1  g478(.A(G8gat), .B1(new_n676), .B2(new_n411), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n676), .A2(new_n411), .A3(new_n682), .ZN(new_n683));
  MUX2_X1   g482(.A(new_n681), .B(KEYINPUT42), .S(new_n683), .Z(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n676), .B2(new_n506), .ZN(new_n685));
  INV_X1    g484(.A(new_n467), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n676), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n676), .A2(new_n293), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n649), .A2(new_n692), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n466), .A2(new_n475), .B1(new_n482), .B2(KEYINPUT35), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n507), .A2(new_n485), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n674), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n607), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n564), .A2(new_n572), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT108), .B1(new_n644), .B2(new_n648), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n634), .A2(new_n636), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT36), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n477), .B(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n282), .A2(new_n292), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n708), .A2(new_n291), .B1(new_n491), .B2(new_n494), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(new_n504), .ZN(new_n710));
  INV_X1    g509(.A(new_n293), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n677), .A2(new_n411), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n481), .B2(new_n293), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n705), .B1(new_n484), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n696), .B(new_n701), .C1(new_n718), .C2(KEYINPUT44), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n677), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n476), .A2(new_n483), .B1(new_n710), .B2(new_n716), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n692), .B1(new_n723), .B2(new_n705), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n724), .A2(KEYINPUT109), .A3(new_n696), .A4(new_n701), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n523), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n727), .B2(new_n726), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n698), .A2(new_n649), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n508), .A2(new_n576), .A3(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n731), .A2(G29gat), .A3(new_n677), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT45), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(G1328gat));
  NOR3_X1   g533(.A1(new_n731), .A2(G36gat), .A3(new_n411), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT46), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n721), .A2(new_n479), .A3(new_n725), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n524), .B2(new_n737), .ZN(G1329gat));
  NOR3_X1   g537(.A1(new_n731), .A2(G43gat), .A3(new_n686), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G43gat), .B1(new_n719), .B2(new_n506), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT47), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n721), .A2(new_n707), .A3(new_n725), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n740), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT111), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n739), .B1(new_n743), .B2(G43gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT47), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n747), .B2(new_n750), .ZN(G1330gat));
  OR3_X1    g550(.A1(new_n731), .A2(G50gat), .A3(new_n293), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n724), .A2(new_n711), .A3(new_n696), .A4(new_n701), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT112), .A2(KEYINPUT48), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n731), .A2(new_n758), .A3(G50gat), .A4(new_n293), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n721), .A2(new_n711), .A3(new_n725), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(G50gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n761), .B2(KEYINPUT48), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(KEYINPUT113), .B(new_n757), .C1(new_n761), .C2(KEYINPUT48), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1331gat));
  INV_X1    g565(.A(new_n723), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n652), .A2(new_n699), .A3(new_n697), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n722), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n479), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n774), .B2(new_n773), .ZN(G1333gat));
  OAI21_X1  g576(.A(G71gat), .B1(new_n769), .B2(new_n506), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n686), .A2(G71gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g580(.A1(new_n770), .A2(new_n711), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n724), .A2(new_n696), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n642), .A2(new_n699), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n674), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n784), .A2(KEYINPUT114), .A3(new_n786), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n722), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n619), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n767), .A2(new_n637), .A3(new_n785), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT51), .Z(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n677), .A2(new_n619), .A3(new_n697), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  NOR3_X1   g595(.A1(new_n697), .A2(G92gat), .A3(new_n411), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G92gat), .B1(new_n787), .B2(new_n411), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n788), .A2(new_n479), .A3(new_n789), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n802), .A2(G92gat), .B1(new_n793), .B2(new_n797), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(G1337gat));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n707), .A3(new_n789), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n686), .A2(G99gat), .A3(new_n697), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n794), .B2(new_n808), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n293), .A2(G106gat), .A3(new_n697), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G106gat), .B1(new_n787), .B2(new_n293), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n788), .A2(new_n711), .A3(new_n789), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n815), .A2(G106gat), .B1(new_n793), .B2(new_n810), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n813), .ZN(G1339gat));
  NAND3_X1  g616(.A1(new_n655), .A2(new_n660), .A3(new_n670), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n668), .B1(new_n671), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n669), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n821), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n823), .B1(new_n822), .B2(new_n669), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n562), .A2(new_n546), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n544), .A2(new_n548), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n513), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n572), .A2(new_n833), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n702), .A2(new_n704), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n822), .A2(new_n669), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n699), .A2(new_n837), .A3(new_n824), .A4(new_n827), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n834), .A2(new_n674), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n702), .A2(new_n704), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n607), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n638), .A2(new_n651), .A3(new_n700), .A4(new_n697), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n677), .A2(new_n479), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n478), .ZN(new_n846));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n699), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n293), .A3(new_n467), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n352), .A3(new_n575), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(G1340gat));
  AOI21_X1  g649(.A(G120gat), .B1(new_n846), .B2(new_n674), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n848), .A2(new_n350), .A3(new_n697), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(G1341gat));
  NAND3_X1  g652(.A1(new_n846), .A2(new_n345), .A3(new_n642), .ZN(new_n854));
  OAI21_X1  g653(.A(G127gat), .B1(new_n848), .B2(new_n607), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1342gat));
  AOI21_X1  g655(.A(new_n677), .B1(new_n841), .B2(new_n842), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n649), .A2(new_n479), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n857), .A2(new_n347), .A3(new_n478), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n848), .B2(new_n649), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  NAND2_X1  g661(.A1(new_n506), .A2(new_n844), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n711), .A2(KEYINPUT57), .ZN(new_n865));
  INV_X1    g664(.A(new_n842), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n836), .B1(new_n826), .B2(new_n825), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(new_n573), .B2(new_n574), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n637), .B1(new_n868), .B2(new_n839), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n607), .B1(new_n869), .B2(new_n835), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n870), .B2(KEYINPUT117), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n607), .C1(new_n869), .C2(new_n835), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n865), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n293), .B1(new_n841), .B2(new_n842), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n864), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877), .B2(new_n575), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n707), .A2(new_n293), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n857), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n575), .A2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(new_n411), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n878), .A2(new_n879), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n699), .B(new_n864), .C1(new_n874), .C2(new_n876), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(G141gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(G141gat), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n881), .A2(G141gat), .A3(new_n479), .A4(new_n575), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g692(.A(new_n877), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n674), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n830), .A2(new_n637), .A3(new_n834), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n607), .B1(new_n869), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n638), .A2(new_n651), .A3(new_n575), .A4(new_n697), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n293), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n674), .A3(new_n864), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n882), .A2(new_n884), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n479), .A3(new_n697), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n895), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n896), .B(new_n907), .C1(new_n910), .C2(G148gat), .ZN(G1345gat));
  NAND4_X1  g710(.A1(new_n882), .A2(new_n411), .A3(new_n642), .A4(new_n884), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n642), .A2(G155gat), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT121), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n912), .A2(new_n232), .B1(new_n894), .B2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n877), .B2(new_n705), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n858), .A2(new_n233), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n916), .B(new_n920), .C1(new_n908), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1347gat));
  NOR3_X1   g721(.A1(new_n394), .A2(new_n722), .A3(new_n411), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n843), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n324), .A3(new_n575), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n843), .A2(new_n677), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n843), .A2(KEYINPUT123), .A3(new_n677), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n478), .A2(new_n479), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n699), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n926), .B1(new_n935), .B2(new_n324), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n925), .B2(new_n697), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n674), .A2(new_n325), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n933), .B2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n925), .B2(new_n607), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n642), .A2(new_n332), .ZN(new_n942));
  OAI221_X1 g741(.A(new_n940), .B1(KEYINPUT124), .B2(new_n941), .C1(new_n933), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(KEYINPUT124), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1350gat));
  OR3_X1    g744(.A1(new_n933), .A2(G190gat), .A3(new_n705), .ZN(new_n946));
  OAI21_X1  g745(.A(G190gat), .B1(new_n925), .B2(new_n649), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT125), .B1(new_n947), .B2(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n947), .A2(KEYINPUT125), .A3(KEYINPUT61), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NAND2_X1  g751(.A1(new_n880), .A2(new_n479), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n931), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n699), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n707), .A2(new_n722), .A3(new_n411), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n905), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n576), .A2(G197gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n959), .B2(new_n697), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n905), .A2(KEYINPUT127), .A3(new_n674), .A4(new_n958), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(G204gat), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n697), .A2(G204gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT123), .B1(new_n843), .B2(new_n677), .ZN(new_n969));
  AOI211_X1 g768(.A(new_n928), .B(new_n722), .C1(new_n841), .C2(new_n842), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n954), .B(new_n968), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n974), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n972), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n966), .A2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n905), .A2(new_n642), .A3(new_n958), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n607), .A2(G211gat), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n981), .A2(new_n982), .B1(new_n955), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n959), .B2(new_n649), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n705), .A2(G218gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n955), .B2(new_n986), .ZN(G1355gat));
endmodule


