//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1185, new_n1186, new_n1187, new_n1188, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G250), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n204), .B1(new_n205), .B2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G13), .ZN(new_n207));
  NAND4_X1  g0007(.A1(new_n207), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n203), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(G20), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n214), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G116), .ZN(new_n224));
  INV_X1    g0024(.A(G270), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  INV_X1    g0029(.A(G97), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n211), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n226), .B(new_n231), .C1(G58), .C2(G232), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(G1), .B2(G20), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT1), .Z(new_n234));
  NOR2_X1   g0034(.A1(new_n222), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n225), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n224), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(G226), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  OAI211_X1 g0055(.A(G232), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G41), .A2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n262), .A2(G1), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT67), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n262), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n259), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G238), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n258), .A2(new_n273), .A3(new_n259), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n261), .A2(new_n265), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n264), .B1(new_n260), .B2(KEYINPUT71), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(new_n272), .A4(new_n274), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(new_n283), .B2(G68), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT72), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  INV_X1    g0088(.A(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n205), .B2(new_n289), .ZN(new_n293));
  NAND4_X1  g0093(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n217), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT11), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT67), .B(G1), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n299), .A2(new_n207), .A3(new_n283), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n228), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n291), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n293), .A2(new_n217), .A3(new_n294), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n283), .B2(new_n299), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G68), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n298), .A2(new_n302), .A3(new_n303), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n276), .B2(new_n279), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n282), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n280), .A2(KEYINPUT73), .A3(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n276), .A2(G179), .A3(new_n279), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n315), .A4(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n311), .B1(new_n317), .B2(new_n308), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT74), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n300), .A2(G50), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(G50), .B2(new_n305), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT69), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  INV_X1    g0123(.A(G150), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n284), .B1(new_n324), .B2(new_n290), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G58), .A2(G68), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n283), .B1(new_n326), .B2(new_n288), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n295), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n271), .A2(G226), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT3), .B(G33), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(G222), .A3(new_n252), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n285), .B2(new_n332), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n289), .ZN(new_n336));
  NAND2_X1  g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n252), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n334), .B1(G223), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G41), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n218), .B1(new_n289), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n265), .B(new_n331), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n342), .A2(G179), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n330), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n329), .A2(KEYINPUT9), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n329), .A2(KEYINPUT9), .B1(G200), .B2(new_n342), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n342), .A2(new_n281), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(KEYINPUT10), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n336), .A2(new_n283), .A3(new_n337), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n283), .A4(new_n337), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n283), .A2(new_n289), .A3(G159), .ZN(new_n361));
  INV_X1    g0161(.A(G58), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n228), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n326), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n360), .A2(KEYINPUT16), .A3(new_n361), .A4(new_n364), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n295), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n306), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n300), .A2(new_n323), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n332), .A2(G226), .A3(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  OAI211_X1 g0175(.A(G223), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n259), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n271), .B2(G232), .ZN(new_n380));
  INV_X1    g0180(.A(G232), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n270), .A2(new_n259), .A3(KEYINPUT75), .A4(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n378), .B(new_n265), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n341), .B1(new_n299), .B2(new_n262), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT75), .B1(new_n389), .B2(new_n381), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n271), .A2(new_n379), .A3(G232), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n392), .A2(KEYINPUT76), .A3(new_n378), .A4(new_n265), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n343), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n373), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n388), .A2(new_n309), .A3(new_n393), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n384), .A2(new_n281), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n373), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n398), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n400), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT77), .B1(new_n399), .B2(new_n400), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n398), .B(new_n406), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n397), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n300), .A2(new_n285), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n306), .A2(G77), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT15), .B(G87), .Z(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n284), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n323), .A2(new_n290), .B1(new_n283), .B2(new_n285), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n295), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n332), .A2(G232), .A3(new_n252), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  INV_X1    g0224(.A(new_n338), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n423), .B1(new_n424), .B2(new_n332), .C1(new_n425), .C2(new_n229), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n259), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n271), .A2(G244), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n265), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n422), .B(new_n430), .C1(new_n281), .C2(new_n429), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n429), .A2(G179), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n343), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n421), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n412), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n319), .A2(new_n354), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n267), .A2(new_n269), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(G13), .A3(G20), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(G33), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n304), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G107), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT85), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n300), .B(new_n424), .C1(new_n445), .C2(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(KEYINPUT25), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n424), .A2(G20), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT84), .B1(new_n449), .B2(KEYINPUT23), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT84), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n424), .A4(G20), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n450), .A2(new_n453), .B1(KEYINPUT23), .B2(new_n449), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n283), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n283), .A2(G33), .A3(G116), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n332), .A2(new_n283), .A3(G87), .A4(new_n458), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n454), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n463), .B(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n444), .B(new_n448), .C1(new_n465), .C2(new_n304), .ZN(new_n466));
  OAI211_X1 g0266(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n467));
  OAI211_X1 g0267(.A(G250), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n468));
  INV_X1    g0268(.A(G294), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(new_n468), .C1(new_n289), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n259), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(KEYINPUT86), .A3(new_n259), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n267), .B2(new_n269), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n259), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G264), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n476), .A2(new_n341), .A3(G274), .A4(new_n477), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n473), .A2(new_n474), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G169), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n471), .A2(new_n479), .A3(new_n480), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n483), .A2(new_n385), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n466), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n309), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n481), .B2(G190), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n463), .B(KEYINPUT24), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n295), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(new_n490), .A3(new_n444), .A4(new_n448), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n332), .A2(G257), .A3(new_n252), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n253), .A2(new_n254), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G303), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n493), .B(new_n495), .C1(new_n425), .C2(new_n212), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n259), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n478), .A2(new_n498), .A3(G270), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n498), .B1(new_n478), .B2(G270), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n480), .B(new_n497), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n224), .A2(G20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n283), .C1(G33), .C2(new_n230), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n295), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n295), .A2(KEYINPUT20), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n300), .A2(new_n224), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n304), .A2(G116), .A3(new_n440), .A4(new_n441), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n502), .A2(G169), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n502), .A2(G200), .ZN(new_n517));
  INV_X1    g0317(.A(new_n480), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n439), .A2(new_n477), .A3(G45), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n341), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT82), .B1(new_n520), .B2(new_n225), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n521), .B2(new_n499), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(G190), .A3(new_n497), .ZN(new_n523));
  INV_X1    g0323(.A(new_n513), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n502), .A2(new_n513), .A3(KEYINPUT21), .A4(G169), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n513), .A2(new_n522), .A3(G179), .A4(new_n497), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n516), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n492), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n230), .A2(new_n424), .A3(KEYINPUT6), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT78), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G97), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n530), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n424), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n532), .A2(G97), .A3(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n230), .A2(KEYINPUT6), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT78), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(G20), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n290), .A2(new_n285), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n359), .B2(G107), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n295), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT79), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT79), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n548), .A3(new_n295), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n519), .A2(G257), .A3(new_n341), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n551), .A2(new_n552), .A3(new_n480), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n551), .B2(new_n480), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n332), .A2(KEYINPUT4), .A3(G244), .A4(new_n252), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n332), .A2(G250), .A3(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n504), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT80), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n338), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT80), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n558), .A4(new_n559), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n341), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(G200), .B1(new_n555), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n259), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n570), .A2(G190), .A3(new_n480), .A4(new_n551), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n440), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n443), .B2(G97), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n550), .A2(new_n568), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n548), .B1(new_n545), .B2(new_n295), .ZN(new_n575));
  AOI211_X1 g0375(.A(KEYINPUT79), .B(new_n304), .C1(new_n542), .C2(new_n544), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n553), .A2(new_n554), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(new_n385), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n551), .A2(new_n480), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n343), .B1(new_n567), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n259), .B1(new_n476), .B2(new_n263), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n203), .B1(new_n299), .B2(new_n475), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G238), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n586));
  OAI211_X1 g0386(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n259), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n585), .A2(new_n590), .A3(G190), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n283), .B1(new_n257), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G87), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n230), .A3(new_n424), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n283), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n592), .B1(new_n257), .B2(G20), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n295), .B1(new_n300), .B2(new_n417), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n304), .A2(G87), .A3(new_n440), .A4(new_n441), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n591), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(new_n590), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n584), .A2(new_n583), .B1(new_n589), .B2(new_n259), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n304), .A2(new_n440), .A3(new_n416), .A4(new_n441), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n606), .A2(new_n385), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n343), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n603), .A2(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n574), .A2(new_n582), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n438), .A2(new_n529), .A3(new_n611), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n352), .A2(new_n353), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT17), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n311), .B1(new_n615), .B2(new_n410), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n317), .A2(new_n308), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n434), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n395), .B(KEYINPUT18), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n613), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n573), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n547), .B2(new_n549), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n579), .A2(new_n581), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  XOR2_X1   g0426(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n627));
  NAND4_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n610), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n590), .A2(KEYINPUT87), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n589), .A2(new_n631), .A3(new_n259), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n632), .B1(new_n584), .B2(new_n583), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n603), .B1(new_n633), .B2(new_n309), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n608), .B1(new_n633), .B2(G169), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n629), .B1(new_n582), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n577), .A2(new_n610), .A3(new_n579), .A4(new_n581), .ZN(new_n638));
  INV_X1    g0438(.A(new_n627), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT89), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n628), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n486), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n516), .A2(new_n526), .A3(new_n527), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n491), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n574), .A2(new_n582), .A3(new_n634), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n635), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n346), .B(new_n621), .C1(new_n437), .C2(new_n647), .ZN(G369));
  NOR2_X1   g0448(.A1(new_n207), .A2(G20), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n299), .A2(new_n650), .A3(KEYINPUT27), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n299), .B2(new_n650), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(G213), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n643), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(new_n492), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n642), .A2(new_n655), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n466), .A2(new_n655), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n486), .A2(new_n660), .A3(new_n491), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n524), .A2(new_n656), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n643), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n528), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n491), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n516), .A2(new_n526), .A3(new_n527), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n486), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n656), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(G399));
  OAI21_X1  g0474(.A(KEYINPUT91), .B1(new_n210), .B2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n210), .A2(KEYINPUT91), .A3(G41), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n595), .A2(G116), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n215), .B2(new_n679), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n656), .B1(new_n641), .B2(new_n646), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT95), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT95), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n688), .B(new_n656), .C1(new_n641), .C2(new_n646), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n582), .A2(new_n636), .A3(new_n629), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n638), .B2(new_n639), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n656), .B1(new_n692), .B2(new_n646), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n567), .A2(new_n580), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n606), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n471), .A2(new_n479), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n522), .A2(G179), .A3(new_n700), .A4(new_n497), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT94), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT93), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n702), .B2(KEYINPUT30), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n698), .A2(new_n701), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n701), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT30), .B1(new_n702), .B2(KEYINPUT93), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n606), .A3(new_n697), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n570), .A2(new_n578), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n633), .A2(G179), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n483), .A4(new_n502), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n656), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g0514(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n696), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n611), .A2(new_n529), .A3(new_n656), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n710), .A2(new_n713), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n655), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(new_n720), .A3(KEYINPUT31), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n695), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n684), .B1(new_n722), .B2(G1), .ZN(G364));
  AOI21_X1  g0523(.A(new_n266), .B1(new_n649), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n678), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n666), .B2(G330), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G330), .B2(new_n666), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n217), .B1(G20), .B2(new_n343), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n283), .A2(G179), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(new_n281), .A3(new_n309), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G329), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n281), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n385), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n734), .B1(new_n738), .B2(new_n469), .ZN(new_n739));
  NAND2_X1  g0539(.A1(G20), .A2(G179), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT97), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n281), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n309), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT33), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(G317), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n745), .B2(G317), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n743), .A2(G200), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n739), .B(new_n747), .C1(G311), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n742), .A2(new_n735), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G322), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n281), .A2(new_n309), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n742), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G326), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n731), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n494), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n752), .B(new_n756), .C1(KEYINPUT98), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(KEYINPUT98), .B2(new_n759), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n731), .A2(new_n281), .A3(G200), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n749), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n332), .B1(new_n757), .B2(new_n594), .C1(new_n424), .C2(new_n763), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n748), .B2(G77), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n744), .A2(G68), .B1(G97), .B2(new_n737), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G50), .A2(new_n755), .B1(new_n751), .B2(G58), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n732), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n730), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n210), .A2(G116), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n729), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n332), .B1(new_n247), .B2(G45), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n216), .A2(new_n475), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n210), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n332), .A2(G355), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n773), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n778), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n666), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n726), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n728), .B1(new_n788), .B2(new_n789), .ZN(G396));
  INV_X1    g0590(.A(new_n635), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n574), .A2(new_n582), .A3(new_n634), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n672), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n628), .A2(new_n640), .A3(new_n637), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n655), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n432), .A2(new_n421), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT100), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n796), .A2(new_n797), .A3(new_n433), .A4(new_n655), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n431), .B(new_n434), .C1(new_n422), .C2(new_n656), .ZN(new_n799));
  OAI21_X1  g0599(.A(KEYINPUT100), .B1(new_n434), .B2(new_n656), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n686), .A2(new_n689), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT102), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n801), .B(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n721), .A2(new_n717), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n806), .B(new_n807), .Z(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n789), .ZN(new_n809));
  INV_X1    g0609(.A(new_n744), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n324), .B1(new_n754), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G159), .B2(new_n748), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n750), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n763), .A2(new_n228), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n332), .B1(new_n732), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(G58), .C2(new_n737), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n816), .B(new_n820), .C1(new_n288), .C2(new_n757), .ZN(new_n821));
  INV_X1    g0621(.A(new_n763), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G87), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n732), .C1(new_n738), .C2(new_n230), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n494), .B1(new_n757), .B2(new_n424), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n758), .B2(new_n754), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G116), .B2(new_n748), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n810), .A2(KEYINPUT99), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n810), .A2(KEYINPUT99), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n829), .B1(new_n762), .B2(new_n832), .C1(new_n469), .C2(new_n750), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n821), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n789), .B1(new_n834), .B2(new_n729), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n729), .A2(new_n775), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(G77), .B2(new_n837), .C1(new_n777), .C2(new_n801), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT101), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n809), .A2(new_n839), .ZN(G384));
  NAND2_X1  g0640(.A1(new_n536), .A2(new_n541), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT35), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n283), .B(new_n217), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(G116), .C1(new_n842), .C2(new_n841), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  OAI21_X1  g0645(.A(G77), .B1(new_n362), .B2(new_n228), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n846), .A2(new_n215), .B1(G50), .B2(new_n228), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n207), .A3(new_n299), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(new_n653), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n373), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n614), .A2(new_n395), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n614), .A2(new_n854), .A3(new_n395), .A4(new_n851), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n615), .A2(new_n410), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n851), .B1(new_n857), .B2(new_n397), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n849), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n851), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n412), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n855), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n718), .A2(new_n720), .A3(new_n715), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT31), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n714), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n801), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n308), .A2(new_n655), .ZN(new_n869));
  INV_X1    g0669(.A(new_n311), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n617), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n869), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n872), .B(new_n311), .C1(new_n317), .C2(new_n308), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n864), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n865), .A2(new_n867), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n437), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n881), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(G330), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n621), .A2(new_n346), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n695), .B2(new_n438), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT104), .Z(new_n888));
  XNOR2_X1  g0688(.A(new_n885), .B(new_n888), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n856), .A2(new_n858), .A3(new_n849), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT39), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n859), .A2(new_n863), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n317), .A2(new_n308), .A3(new_n656), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n620), .A2(new_n653), .ZN(new_n899));
  INV_X1    g0699(.A(new_n874), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n434), .A2(new_n655), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n795), .B2(new_n801), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n864), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n898), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n889), .B(new_n905), .Z(new_n906));
  NOR2_X1   g0706(.A1(new_n439), .A2(new_n649), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n845), .B(new_n848), .C1(new_n906), .C2(new_n907), .ZN(G367));
  INV_X1    g0708(.A(new_n748), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n832), .A2(new_n769), .B1(new_n288), .B2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n910), .A2(KEYINPUT110), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n737), .A2(G68), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(KEYINPUT110), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n811), .A2(new_n732), .B1(new_n757), .B2(new_n362), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT112), .Z(new_n915));
  OAI21_X1  g0715(.A(new_n332), .B1(new_n763), .B2(new_n285), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT111), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n814), .A2(new_n754), .B1(new_n750), .B2(new_n324), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n919), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n494), .B1(new_n750), .B2(new_n758), .C1(new_n824), .C2(new_n754), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(G317), .B2(new_n733), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n763), .A2(new_n230), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G107), .B2(new_n737), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n909), .B2(new_n762), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n922), .B(new_n926), .C1(new_n832), .C2(new_n469), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n757), .A2(new_n224), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT46), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n789), .B1(new_n932), .B2(new_n729), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n209), .A2(new_n494), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n779), .B1(new_n209), .B2(new_n417), .C1(new_n243), .C2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n655), .A2(new_n602), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n634), .A2(new_n635), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(new_n635), .C2(new_n937), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n933), .B(new_n936), .C1(new_n787), .C2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n678), .B(KEYINPUT41), .Z(new_n943));
  XOR2_X1   g0743(.A(new_n663), .B(new_n667), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n722), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n574), .A2(new_n582), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n623), .B2(new_n656), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n625), .A2(new_n655), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n673), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT107), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n950), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n673), .A2(new_n946), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT44), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n953), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n945), .A2(KEYINPUT108), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n943), .B1(new_n960), .B2(new_n722), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n725), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n582), .B1(new_n947), .B2(new_n486), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT106), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(new_n655), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n947), .A2(new_n658), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT42), .Z(new_n968));
  OAI21_X1  g0768(.A(new_n963), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n668), .A2(new_n949), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n942), .B1(new_n962), .B2(new_n973), .ZN(G387));
  OR2_X1    g0774(.A1(new_n722), .A2(new_n944), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT115), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n977), .A2(new_n678), .A3(new_n945), .A4(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n733), .A2(G326), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n909), .A2(new_n758), .B1(new_n750), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n832), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(G311), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT114), .B(G322), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n754), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT48), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n762), .B2(new_n738), .C1(new_n469), .C2(new_n757), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT49), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n332), .B(new_n980), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n989), .B2(new_n988), .C1(new_n224), .C2(new_n763), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n737), .A2(new_n416), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n285), .B2(new_n757), .C1(new_n324), .C2(new_n732), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n288), .A2(new_n750), .B1(new_n754), .B2(new_n769), .ZN(new_n994));
  NOR4_X1   g0794(.A1(new_n993), .A2(new_n994), .A3(new_n494), .A4(new_n923), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n228), .B2(new_n909), .C1(new_n323), .C2(new_n810), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n730), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n370), .A2(new_n288), .ZN(new_n998));
  AOI21_X1  g0798(.A(G45), .B1(new_n998), .B2(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(KEYINPUT50), .B2(new_n998), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G68), .B2(G77), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n681), .B1(new_n1001), .B2(new_n332), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n240), .A2(G45), .A3(new_n494), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n210), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n780), .B(new_n1004), .C1(G107), .C2(new_n210), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n659), .A2(new_n661), .A3(new_n778), .ZN(new_n1006));
  OR4_X1    g0806(.A1(new_n789), .A2(new_n997), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n944), .A2(new_n725), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n979), .A2(new_n1007), .A3(new_n1008), .ZN(G393));
  OAI22_X1  g0809(.A1(new_n832), .A2(new_n758), .B1(new_n224), .B2(new_n738), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT118), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n494), .B1(new_n762), .B2(new_n757), .C1(new_n909), .C2(new_n469), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n824), .A2(new_n750), .B1(new_n754), .B2(new_n981), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT117), .Z(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1014), .B2(KEYINPUT52), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n985), .A2(new_n732), .B1(new_n763), .B2(new_n424), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1011), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n983), .A2(G50), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G150), .A2(new_n755), .B1(new_n751), .B2(G159), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT51), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G143), .A2(new_n733), .B1(new_n737), .B2(G77), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n228), .B2(new_n757), .C1(new_n909), .C2(new_n323), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1021), .A2(KEYINPUT51), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1020), .A2(new_n1026), .A3(new_n332), .A4(new_n823), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1019), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n789), .B1(new_n1028), .B2(new_n729), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n779), .B1(new_n230), .B2(new_n209), .C1(new_n250), .C2(new_n934), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT116), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(new_n787), .C2(new_n949), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n959), .B(new_n669), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n679), .B1(new_n1034), .B2(new_n945), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1033), .B1(new_n1035), .B2(new_n960), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n724), .B2(new_n1034), .ZN(G390));
  NOR3_X1   g0837(.A1(new_n868), .A2(new_n874), .A3(new_n696), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n721), .A2(new_n717), .A3(new_n801), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(new_n874), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n903), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n805), .A2(G330), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n874), .B1(new_n1042), .B2(new_n882), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1039), .A2(new_n874), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n656), .B(new_n801), .C1(new_n692), .C2(new_n646), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n901), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n883), .A2(G330), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n887), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n896), .B1(new_n902), .B2(new_n874), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n892), .A2(new_n894), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n864), .B(new_n896), .C1(new_n874), .C2(new_n1047), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1038), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1044), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1051), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT119), .B1(new_n1060), .B2(new_n679), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1038), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n1051), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT119), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n678), .C1(new_n1064), .C2(new_n1051), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1061), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(KEYINPUT120), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT120), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1061), .A2(new_n1067), .A3(new_n1070), .A4(new_n1065), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n983), .A2(G137), .B1(G159), .B2(new_n737), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT54), .B(G143), .Z(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n909), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT121), .Z(new_n1077));
  INV_X1    g0877(.A(G125), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n332), .B1(new_n763), .B2(new_n288), .C1(new_n1078), .C2(new_n732), .ZN(new_n1079));
  INV_X1    g0879(.A(G128), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1080), .A2(new_n754), .B1(new_n750), .B2(new_n818), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n757), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(G150), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .A4(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n494), .B1(new_n230), .B2(new_n909), .C1(new_n832), .C2(new_n424), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n224), .A2(new_n750), .B1(new_n754), .B2(new_n762), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G294), .A2(new_n733), .B1(new_n737), .B2(G77), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n594), .B2(new_n757), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1086), .A2(new_n817), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n789), .B1(new_n1091), .B2(new_n729), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n370), .B2(new_n837), .C1(new_n895), .C2(new_n777), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1064), .B2(new_n724), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1072), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT122), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT122), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1072), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(G378));
  INV_X1    g0900(.A(new_n1049), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n887), .B(new_n1050), .C1(new_n1064), .C2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n878), .A2(G330), .A3(new_n879), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n905), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n329), .A2(new_n653), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n354), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n354), .A2(new_n1106), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT55), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n354), .A2(new_n1106), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT55), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n1107), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT56), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n878), .A2(G330), .A3(new_n879), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1116), .A2(new_n899), .A3(new_n898), .A4(new_n904), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1104), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1104), .B2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1102), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(KEYINPUT57), .B(new_n1102), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n678), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1115), .A2(new_n776), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n755), .A2(G125), .B1(G150), .B2(new_n737), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1080), .B2(new_n750), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n818), .A2(new_n810), .B1(new_n909), .B2(new_n811), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n1082), .C2(new_n1074), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT59), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G41), .B1(new_n733), .B2(G124), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G33), .B1(new_n822), .B2(G159), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n340), .B(new_n494), .C1(new_n757), .C2(new_n285), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n822), .A2(G58), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1135), .B(new_n912), .C1(new_n762), .C2(new_n732), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G107), .C2(new_n751), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G97), .A2(new_n744), .B1(new_n748), .B2(new_n416), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n224), .C2(new_n754), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT58), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n288), .B1(new_n253), .B2(G41), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1133), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT123), .Z(new_n1143));
  AOI21_X1  g0943(.A(new_n789), .B1(new_n1143), .B2(new_n729), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1125), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n288), .B2(new_n836), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n725), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1124), .A2(new_n1148), .ZN(G375));
  NAND2_X1  g0949(.A1(new_n887), .A2(new_n1050), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1101), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT124), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1101), .A3(KEYINPUT124), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n943), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n1051), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1049), .A2(new_n725), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n874), .A2(new_n775), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n992), .B1(new_n285), .B2(new_n763), .C1(new_n758), .C2(new_n732), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n494), .B1(new_n757), .B2(new_n230), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n469), .B2(new_n754), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n832), .A2(new_n224), .B1(new_n424), .B2(new_n909), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT125), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n1165), .B2(new_n1164), .C1(new_n762), .C2(new_n750), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1135), .B1(new_n750), .B2(new_n811), .C1(new_n818), .C2(new_n754), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G150), .B2(new_n748), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n738), .A2(new_n288), .B1(new_n732), .B2(new_n1080), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n494), .B(new_n1170), .C1(G159), .C2(new_n1082), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n832), .C2(new_n1075), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n789), .B1(new_n1173), .B2(new_n729), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1159), .B(new_n1174), .C1(G68), .C2(new_n837), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1157), .A2(new_n1158), .A3(new_n1175), .ZN(G381));
  NOR2_X1   g0976(.A1(new_n1034), .A2(new_n724), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1033), .B(new_n1177), .C1(new_n960), .C2(new_n1035), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n942), .C1(new_n962), .C2(new_n973), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1179), .A2(G396), .A3(G393), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1068), .A2(new_n1095), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(G375), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G381), .A2(G384), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(G407));
  NAND2_X1  g0984(.A1(new_n654), .A2(G213), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT126), .Z(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(G407), .A2(G213), .A3(new_n1188), .ZN(G409));
  NAND2_X1  g0989(.A1(G387), .A2(G390), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1179), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(G393), .B(G396), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1191), .B(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1158), .A2(new_n1175), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT60), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1151), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1051), .A2(KEYINPUT60), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1155), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1199), .B2(new_n678), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT127), .B1(new_n1200), .B2(G384), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(G384), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT127), .ZN(new_n1203));
  INV_X1    g1003(.A(G384), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n679), .B(new_n1197), .C1(new_n1155), .C2(new_n1198), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1204), .C1(new_n1205), .C2(new_n1195), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G375), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1147), .A2(new_n1156), .A3(new_n1102), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1181), .B1(new_n1148), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1185), .B(new_n1208), .C1(new_n1209), .C2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT62), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1124), .A2(new_n1148), .ZN(new_n1214));
  AOI211_X1 g1014(.A(KEYINPUT122), .B(new_n1094), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1098), .B1(new_n1072), .B2(new_n1095), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1211), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1187), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1212), .A2(new_n1213), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1207), .A2(G2897), .A3(new_n1187), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n654), .A2(G213), .A3(G2897), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1201), .A2(new_n1224), .A3(new_n1202), .A4(new_n1206), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1222), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1194), .B1(new_n1221), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1207), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1194), .B1(new_n1219), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1185), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1226), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1212), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1222), .B(new_n1231), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1228), .A2(new_n1236), .ZN(G405));
  NOR2_X1   g1037(.A1(new_n1214), .A2(new_n1181), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1194), .A2(new_n1217), .A3(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1191), .B(new_n1192), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1238), .B2(new_n1209), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1207), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1242), .A3(new_n1208), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(G402));
endmodule


