//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  MUX2_X1   g049(.A(G100), .B(G112), .S(G2105), .Z(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G124), .B1(G2104), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  INV_X1    g052(.A(new_n463), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT67), .Z(G162));
  INV_X1    g055(.A(G126), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n483), .B2(new_n484), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n489), .C1(new_n460), .C2(new_n461), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G50), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n501), .A2(KEYINPUT6), .A3(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT6), .B1(new_n501), .B2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n500), .A2(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n510), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n510), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n502), .A2(new_n503), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n522), .A2(new_n507), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n520), .A2(new_n524), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT71), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n515), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n505), .B1(new_n511), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n523), .A2(G81), .B1(new_n525), .B2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(KEYINPUT72), .B(new_n538), .C1(new_n541), .C2(new_n515), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n515), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  INV_X1    g119(.A(new_n538), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n521), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(KEYINPUT74), .A3(G651), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n559), .A2(new_n560), .B1(G91), .B2(new_n523), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n505), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n525), .A2(new_n564), .A3(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT73), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n561), .A2(new_n567), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  OR2_X1    g146(.A1(new_n513), .A2(new_n516), .ZN(G303));
  OAI21_X1  g147(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n523), .A2(G87), .B1(new_n525), .B2(G49), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n504), .A2(G86), .A3(new_n510), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(new_n577), .B1(new_n525), .B2(G48), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n508), .B2(new_n509), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT75), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n523), .A2(KEYINPUT76), .A3(G86), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n578), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n515), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT77), .B(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n523), .A2(G85), .B1(new_n525), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT78), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n521), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n525), .B2(G54), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n511), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G168), .B2(new_n610), .ZN(G297));
  XOR2_X1   g187(.A(G297), .B(KEYINPUT80), .Z(G280));
  XNOR2_X1  g188(.A(KEYINPUT81), .B(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(G860), .B2(new_n614), .ZN(G148));
  NAND2_X1  g190(.A1(new_n547), .A2(new_n610), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n604), .A2(new_n605), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n600), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT79), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n606), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n619), .A2(new_n621), .A3(new_n614), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(new_n610), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n463), .A2(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n627), .A2(KEYINPUT13), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(KEYINPUT13), .B2(new_n627), .ZN(new_n631));
  OR3_X1    g206(.A1(new_n631), .A2(new_n628), .A3(new_n629), .ZN(new_n632));
  MUX2_X1   g207(.A(G99), .B(G111), .S(G2105), .Z(new_n633));
  AOI22_X1  g208(.A1(new_n474), .A2(G123), .B1(G2104), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n478), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n631), .B1(new_n628), .B2(new_n629), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n632), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT86), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n667), .B2(new_n661), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n661), .B(KEYINPUT17), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n669), .B(new_n670), .C1(new_n667), .C2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n667), .A3(new_n664), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n629), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT89), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  OR2_X1    g260(.A1(new_n678), .A2(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n683), .A3(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n683), .C2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(G229));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n695), .B(new_n697), .Z(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G22), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G166), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n698), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n710));
  MUX2_X1   g285(.A(G24), .B(G290), .S(G16), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(G1986), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(G1986), .ZN(new_n713));
  MUX2_X1   g288(.A(G95), .B(G107), .S(G2105), .Z(new_n714));
  AOI22_X1  g289(.A1(new_n474), .A2(G119), .B1(G2104), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G131), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n478), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT90), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n710), .A2(new_n712), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n726), .A2(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n726), .A2(KEYINPUT92), .A3(KEYINPUT36), .A4(new_n727), .ZN(new_n732));
  NOR2_X1   g307(.A1(G29), .A2(G33), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT25), .B1(new_n465), .B2(G103), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n489), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n736), .B(new_n738), .C1(G139), .C2(new_n463), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n719), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n719), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n743), .B1(G2090), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n699), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n547), .B2(new_n699), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n699), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n699), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1961), .ZN(new_n753));
  INV_X1    g328(.A(new_n746), .ZN(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n747), .A2(new_n750), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n699), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n699), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1966), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n741), .A2(G2072), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n699), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n607), .B2(new_n699), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT93), .B(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n699), .A2(G20), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  INV_X1    g344(.A(G299), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n699), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1956), .Z(new_n772));
  OR2_X1    g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  NAND2_X1  g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G160), .B2(G29), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n637), .A2(G29), .B1(new_n776), .B2(G2084), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT26), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G105), .B2(new_n465), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n463), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n474), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n719), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n719), .B2(G32), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n777), .B1(G2084), .B2(new_n776), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT30), .B(G28), .Z(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G29), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n786), .B2(new_n787), .ZN(new_n792));
  NAND2_X1  g367(.A1(G164), .A2(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G27), .B2(G29), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n719), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n474), .A2(G128), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n463), .A2(G140), .ZN(new_n801));
  MUX2_X1   g376(.A(G104), .B(G116), .S(G2105), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G2104), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n719), .ZN(new_n806));
  INV_X1    g381(.A(G2067), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n792), .A2(new_n796), .A3(new_n797), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n788), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n763), .A2(new_n767), .A3(new_n772), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n757), .A2(new_n761), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n731), .A2(new_n732), .A3(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  INV_X1    g389(.A(G55), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n815), .A2(new_n505), .B1(new_n511), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n515), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n607), .A2(G559), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n547), .B1(new_n822), .B2(new_n820), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n823), .B1(new_n544), .B2(new_n545), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n829), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n836), .B(new_n824), .C1(KEYINPUT100), .C2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(KEYINPUT100), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(G162), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n637), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n717), .B(KEYINPUT101), .Z(new_n843));
  MUX2_X1   g418(.A(G106), .B(G118), .S(G2105), .Z(new_n844));
  AOI22_X1  g419(.A1(new_n474), .A2(G130), .B1(G2104), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G142), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n478), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n627), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT102), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n739), .B(new_n784), .ZN(new_n851));
  XNOR2_X1  g426(.A(G164), .B(new_n804), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n854), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n842), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n850), .A2(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n854), .A2(new_n849), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n842), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT40), .Z(G395));
  NOR3_X1   g439(.A1(new_n820), .A2(G868), .A3(new_n822), .ZN(new_n865));
  XNOR2_X1  g440(.A(G290), .B(G288), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(G305), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n866), .B(new_n867), .Z(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n607), .B2(new_n614), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n619), .A2(KEYINPUT103), .A3(new_n621), .A4(new_n614), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n832), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n876), .A2(new_n831), .A3(new_n830), .A4(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n618), .A2(G299), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n606), .A2(new_n561), .A3(new_n567), .A4(new_n569), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n874), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n878), .B2(new_n880), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n878), .A2(new_n880), .A3(new_n884), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(KEYINPUT104), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n874), .A2(new_n877), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n883), .B1(KEYINPUT105), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n874), .A2(new_n877), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n888), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT105), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n870), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n874), .A2(new_n877), .A3(new_n882), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n898), .A2(KEYINPUT42), .A3(new_n893), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n869), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n890), .A2(new_n894), .A3(new_n870), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT42), .B1(new_n898), .B2(new_n893), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n868), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n865), .B1(new_n904), .B2(G868), .ZN(G295));
  AOI21_X1  g480(.A(new_n865), .B1(new_n904), .B2(G868), .ZN(G331));
  XNOR2_X1  g481(.A(G286), .B(G171), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n832), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n832), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n882), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n885), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n908), .A2(new_n909), .B1(new_n886), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n868), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n892), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n869), .A3(new_n910), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n917), .A3(new_n858), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n910), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n868), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n858), .A4(new_n917), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n922), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(KEYINPUT43), .A3(new_n858), .A4(new_n917), .ZN(new_n926));
  XOR2_X1   g501(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(G397));
  NOR2_X1   g504(.A1(G290), .A2(G1986), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n804), .B(new_n807), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n783), .A2(G1996), .ZN(new_n933));
  INV_X1    g508(.A(G1996), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n784), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n723), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n717), .B(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n931), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n498), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  AND4_X1   g525(.A1(KEYINPUT110), .A2(new_n498), .A3(new_n950), .A4(new_n944), .ZN(new_n951));
  AND2_X1   g526(.A1(KEYINPUT4), .A2(G138), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n460), .B2(new_n461), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n492), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n954), .A2(new_n489), .B1(new_n496), .B2(new_n495), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n955), .B2(new_n488), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT110), .B1(new_n956), .B2(new_n950), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n950), .B1(new_n498), .B2(new_n944), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n951), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n943), .ZN(new_n961));
  INV_X1    g536(.A(G2084), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n947), .A2(new_n942), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1966), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G8), .ZN(new_n969));
  NAND2_X1  g544(.A1(G286), .A2(G8), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(KEYINPUT124), .A3(KEYINPUT51), .A4(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n963), .B2(new_n967), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(G286), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n970), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT51), .B1(new_n973), .B2(KEYINPUT124), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n956), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n964), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n980), .A2(new_n982), .A3(new_n942), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n947), .A2(KEYINPUT107), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n945), .A2(new_n985), .A3(new_n946), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n707), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n989), .A2(new_n990), .B1(new_n755), .B2(new_n961), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(KEYINPUT109), .A3(new_n707), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n972), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G166), .A2(new_n972), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT112), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT111), .B(new_n997), .C1(G166), .C2(new_n972), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT55), .B1(new_n994), .B2(new_n995), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n493), .B1(new_n472), .B2(new_n952), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n497), .B1(new_n1003), .B2(G2105), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n472), .A2(G126), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n489), .B1(new_n1005), .B2(new_n486), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n950), .B(new_n944), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n959), .A2(new_n942), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n755), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n972), .B1(new_n989), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n942), .A2(new_n956), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1012), .B(G8), .C1(new_n1013), .C2(G288), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT113), .B(G1976), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(G288), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1012), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(G48), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n576), .B1(new_n505), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G1981), .B1(new_n1022), .B2(new_n584), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G305), .B2(G1981), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT49), .B(new_n1023), .C1(G305), .C2(G1981), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT114), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1019), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1002), .A2(new_n1011), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n980), .A2(new_n982), .A3(new_n942), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n984), .B2(new_n986), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n795), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n466), .A2(KEYINPUT53), .A3(G40), .A4(new_n795), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n469), .B(KEYINPUT125), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(G2105), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1043), .A2(new_n947), .A3(new_n982), .A4(new_n980), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n960), .B2(new_n943), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n956), .A2(KEYINPUT110), .A3(new_n950), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1007), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1050), .B2(new_n958), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(KEYINPUT118), .A3(new_n942), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G1961), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1045), .A2(G171), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1054), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n965), .A2(new_n1039), .A3(G2078), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1035), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(G171), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(G301), .A3(new_n1058), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(KEYINPUT54), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n979), .A2(new_n1034), .A3(new_n1060), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n542), .A2(new_n546), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n983), .A2(new_n987), .A3(new_n934), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1012), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(KEYINPUT121), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1069), .B(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n563), .B2(new_n565), .ZN(new_n1073));
  AOI22_X1  g648(.A1(G299), .A2(KEYINPUT57), .B1(new_n561), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1008), .A2(G1956), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n983), .A2(new_n987), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT117), .B1(new_n1037), .B2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1037), .A2(KEYINPUT117), .A3(new_n1077), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1072), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1075), .B(KEYINPUT120), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(KEYINPUT61), .A3(new_n1085), .A4(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1012), .A2(G2067), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1051), .A2(KEYINPUT118), .A3(new_n942), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT118), .B1(new_n1051), .B2(new_n942), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1348), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1047), .A2(new_n1099), .A3(new_n1052), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1095), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n606), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1094), .B(new_n1101), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1100), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n618), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1094), .B1(new_n1114), .B2(new_n1101), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1093), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  OR3_X1    g691(.A1(new_n1100), .A2(KEYINPUT119), .A3(new_n618), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n1100), .B2(new_n618), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1090), .A3(new_n1091), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1085), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1064), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1013), .B(new_n701), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G305), .A2(G1981), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT115), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1020), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n972), .B(G286), .C1(new_n963), .C2(new_n967), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(new_n1127), .C1(new_n1001), .C2(new_n1010), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1002), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1129), .B2(new_n1033), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n991), .A2(new_n992), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1033), .A3(new_n1126), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n993), .A2(KEYINPUT116), .A3(new_n1001), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT63), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  AND4_X1   g711(.A1(new_n1059), .A2(new_n1002), .A3(new_n1011), .A4(new_n1033), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT62), .B1(new_n975), .B2(new_n978), .ZN(new_n1138));
  AND4_X1   g713(.A1(KEYINPUT62), .A2(new_n978), .A3(new_n971), .A4(new_n974), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n949), .B1(new_n1121), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n948), .A2(new_n934), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT46), .Z(new_n1144));
  INV_X1    g719(.A(new_n948), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n784), .B2(new_n932), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT47), .Z(new_n1148));
  OR2_X1    g723(.A1(new_n717), .A2(new_n937), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n936), .A2(new_n1149), .B1(G2067), .B2(new_n804), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n948), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n939), .A2(new_n1145), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n931), .A2(new_n1145), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1148), .A2(new_n1151), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1142), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g734(.A1(G229), .A2(new_n458), .A3(G227), .ZN(new_n1161));
  NOR3_X1   g735(.A1(new_n863), .A2(G401), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g736(.A1(new_n1162), .A2(new_n926), .A3(new_n925), .ZN(G308));
  NAND3_X1  g737(.A1(new_n1162), .A2(new_n925), .A3(new_n926), .ZN(G225));
endmodule


