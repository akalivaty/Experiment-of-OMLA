//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(new_n205), .B2(new_n206), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT28), .B1(new_n212), .B2(new_n213), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n209), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n222), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n232), .A3(new_n207), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT25), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT25), .A4(new_n207), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(new_n224), .B2(new_n222), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT65), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n213), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n233), .B(KEYINPUT25), .C1(new_n226), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n230), .A2(new_n232), .A3(new_n207), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n227), .B1(new_n209), .B2(new_n223), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n246), .B2(new_n228), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n242), .B(new_n243), .C1(new_n247), .C2(KEYINPUT25), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n219), .B1(new_n237), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G127gat), .ZN(new_n251));
  INV_X1    g050(.A(G127gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G134gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G120gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G113gat), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n264), .A3(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n249), .A2(new_n269), .ZN(new_n272));
  INV_X1    g071(.A(G227gat), .ZN(new_n273));
  INV_X1    g072(.A(G233gat), .ZN(new_n274));
  OAI22_X1  g073(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT34), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  OAI221_X1 g076(.A(new_n277), .B1(new_n273), .B2(new_n274), .C1(new_n271), .C2(new_n272), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n239), .B(new_n240), .C1(new_n226), .C2(new_n227), .ZN(new_n282));
  INV_X1    g081(.A(new_n228), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n281), .B1(new_n284), .B2(new_n244), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n243), .B1(new_n285), .B2(new_n242), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT65), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n218), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n269), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n274), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n270), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G43gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n293), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n292), .B2(KEYINPUT32), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(KEYINPUT67), .A3(new_n295), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n292), .B(KEYINPUT32), .C1(new_n294), .C2(new_n298), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n280), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n279), .B(new_n308), .C1(new_n302), .C2(new_n304), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n202), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n303), .A2(KEYINPUT67), .A3(new_n295), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT67), .B1(new_n303), .B2(new_n295), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n279), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n280), .B(new_n306), .C1(new_n311), .C2(new_n312), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(KEYINPUT36), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G22gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G155gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT73), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT72), .B(G155gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n328), .B(KEYINPUT2), .C1(new_n329), .C2(new_n320), .ZN(new_n330));
  XOR2_X1   g129(.A(G155gat), .B(G162gat), .Z(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n336), .ZN(new_n340));
  XOR2_X1   g139(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G211gat), .B(G218gat), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n351), .A2(new_n352), .B1(G211gat), .B2(G218gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n351), .B2(new_n352), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT78), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI211_X1 g159(.A(KEYINPUT29), .B(new_n357), .C1(new_n360), .C2(KEYINPUT78), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n348), .B1(new_n361), .B2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n358), .B2(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n355), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n349), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT69), .A3(new_n356), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(KEYINPUT29), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n360), .B2(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n344), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(G228gat), .A3(G233gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT31), .B(G50gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n372), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n372), .B2(new_n377), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n319), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n372), .A2(new_n377), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n372), .A2(new_n377), .A3(new_n379), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n318), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n338), .A2(new_n343), .A3(new_n264), .A4(new_n256), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n256), .A2(new_n264), .A3(KEYINPUT74), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT74), .B1(new_n256), .B2(new_n264), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n339), .A2(new_n334), .A3(new_n335), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT2), .B1(new_n329), .B2(new_n320), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(KEYINPUT73), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n342), .B1(new_n397), .B2(new_n330), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n398), .B2(new_n373), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n388), .B(new_n391), .C1(new_n399), .C2(new_n370), .ZN(new_n400));
  INV_X1    g199(.A(new_n347), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n346), .B1(new_n338), .B2(new_n343), .ZN(new_n402));
  NOR4_X1   g201(.A1(new_n401), .A2(new_n402), .A3(new_n269), .A4(new_n390), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT76), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n388), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n373), .B1(new_n338), .B2(new_n343), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n265), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n256), .A2(new_n264), .A3(KEYINPUT74), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n398), .A2(new_n373), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n345), .A2(new_n289), .A3(KEYINPUT4), .A4(new_n347), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .A4(new_n391), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n389), .B1(new_n410), .B2(new_n398), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND4_X1  g224(.A1(new_n345), .A2(new_n289), .A3(new_n390), .A4(new_n347), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n413), .A3(new_n418), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  INV_X1    g231(.A(new_n420), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n404), .B2(new_n416), .ZN(new_n434));
  INV_X1    g233(.A(new_n429), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT6), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n218), .B(new_n440), .C1(new_n286), .C2(new_n287), .ZN(new_n441));
  INV_X1    g240(.A(new_n369), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n218), .B1(new_n234), .B2(new_n236), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n440), .A2(KEYINPUT29), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n218), .B(new_n440), .C1(new_n234), .C2(new_n236), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n288), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT70), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT30), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(KEYINPUT70), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n444), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n447), .B1(new_n249), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n369), .ZN(new_n461));
  INV_X1    g260(.A(new_n453), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n446), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n456), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n439), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n310), .A2(new_n316), .B1(new_n387), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n411), .A2(new_n412), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n428), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n405), .ZN(new_n471));
  INV_X1    g270(.A(new_n419), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(new_n388), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n426), .A2(new_n427), .B1(new_n412), .B2(new_n411), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n388), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n475), .A3(new_n425), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n471), .A2(new_n475), .A3(KEYINPUT40), .A4(new_n425), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n478), .A2(new_n436), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n387), .B1(new_n480), .B2(new_n464), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n450), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n482), .B1(new_n449), .B2(new_n442), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n441), .A2(new_n445), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n369), .ZN(new_n490));
  AOI211_X1 g289(.A(KEYINPUT38), .B(new_n453), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n487), .A2(new_n491), .B1(new_n450), .B2(new_n453), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n461), .A2(KEYINPUT37), .A3(new_n446), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(new_n462), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n484), .B(KEYINPUT37), .C1(new_n461), .C2(new_n446), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT79), .B1(new_n450), .B2(new_n482), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT38), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(new_n438), .A3(new_n498), .A4(new_n437), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n307), .A2(new_n309), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n382), .A2(new_n386), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n464), .B1(new_n438), .B2(new_n437), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n314), .A2(new_n503), .A3(new_n315), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT35), .B1(new_n506), .B2(new_n466), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n467), .A2(new_n500), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT14), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n511), .B(new_n513), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  INV_X1    g313(.A(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G43gat), .ZN(new_n516));
  INV_X1    g315(.A(G43gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G50gat), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT15), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(KEYINPUT81), .A3(G50gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT80), .B(KEYINPUT15), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n518), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n514), .A2(new_n519), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT17), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(new_n530), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G8gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(G1gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n541), .B2(G1gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n538), .A3(new_n542), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT84), .Z(new_n548));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n549));
  INV_X1    g348(.A(new_n545), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n543), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n544), .A2(KEYINPUT85), .A3(new_n545), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n528), .A2(new_n530), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n546), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n548), .B(KEYINPUT13), .Z(new_n560));
  NOR2_X1   g359(.A1(new_n553), .A2(new_n531), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT86), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT86), .B(new_n560), .C1(new_n556), .C2(new_n561), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n558), .A2(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT11), .B(G169gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n546), .A2(new_n557), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT18), .A3(new_n548), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n572), .B1(new_n566), .B2(new_n574), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT87), .B1(new_n508), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n505), .A2(new_n507), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n466), .A2(new_n387), .ZN(new_n582));
  INV_X1    g381(.A(new_n316), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT36), .B1(new_n314), .B2(new_n315), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n500), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G218gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT8), .ZN(new_n595));
  AND2_X1   g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  OAI221_X1 g395(.A(new_n594), .B1(G85gat), .B2(G92gat), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(G85gat), .B(G92gat), .C1(KEYINPUT92), .C2(KEYINPUT7), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(KEYINPUT92), .B2(KEYINPUT7), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT93), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(KEYINPUT93), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT93), .B(new_n601), .C1(new_n597), .C2(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(KEYINPUT94), .A3(new_n605), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n536), .B2(new_n533), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(new_n555), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n611), .A2(G190gat), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n537), .A2(new_n614), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n213), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n590), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n621));
  OAI21_X1  g420(.A(G190gat), .B1(new_n611), .B2(new_n615), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n618), .A3(new_n213), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(G218gat), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n623), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT91), .B1(new_n628), .B2(new_n590), .ZN(new_n629));
  INV_X1    g428(.A(new_n626), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n630), .A3(new_n624), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  XOR2_X1   g436(.A(G57gat), .B(G64gat), .Z(new_n638));
  AOI211_X1 g437(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(KEYINPUT9), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(KEYINPUT9), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT88), .B(G57gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(G64gat), .ZN(new_n642));
  INV_X1    g441(.A(G64gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(G57gat), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n252), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n554), .B1(new_n648), .B2(new_n647), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT89), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G155gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G183gat), .B(G211gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT90), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n627), .A2(new_n631), .A3(new_n633), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n646), .A4(new_n609), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT95), .B1(new_n597), .B2(new_n599), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(new_n601), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n601), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n647), .A2(new_n604), .A3(new_n605), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n666), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n666), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  OR2_X1    g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n667), .A2(new_n674), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n665), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n666), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n680), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n635), .A2(new_n663), .A3(new_n664), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n589), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT97), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n589), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n439), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  AND3_X1   g497(.A1(new_n694), .A2(new_n464), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n538), .B1(new_n694), .B2(new_n464), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT42), .B2(new_n699), .ZN(G1325gat));
  INV_X1    g501(.A(G15gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n694), .A2(new_n703), .A3(new_n501), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n310), .A2(new_n316), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n691), .B2(new_n693), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(new_n703), .ZN(G1326gat));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n694), .B2(new_n387), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AOI211_X1 g509(.A(KEYINPUT98), .B(new_n503), .C1(new_n691), .C2(new_n693), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n713), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n709), .B2(new_n711), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1327gat));
  NAND2_X1  g516(.A1(new_n635), .A2(new_n664), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n508), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n508), .B2(new_n719), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n579), .A2(new_n663), .A3(new_n686), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n439), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n663), .A2(new_n686), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n580), .B2(new_n588), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n509), .A3(new_n695), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n727), .A2(new_n733), .A3(new_n734), .ZN(G1328gat));
  OAI21_X1  g534(.A(G36gat), .B1(new_n726), .B2(new_n465), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n730), .A2(new_n510), .A3(new_n464), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(KEYINPUT99), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(KEYINPUT99), .ZN(new_n740));
  OAI221_X1 g539(.A(new_n736), .B1(KEYINPUT46), .B2(new_n737), .C1(new_n739), .C2(new_n740), .ZN(G1329gat));
  INV_X1    g540(.A(new_n705), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n742), .A3(new_n723), .A4(new_n725), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n517), .A3(new_n501), .A4(new_n728), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT100), .B1(new_n589), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT100), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n748), .B(new_n745), .C1(new_n580), .C2(new_n588), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n744), .B(KEYINPUT47), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n747), .B2(new_n749), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n587), .B1(new_n586), .B2(new_n578), .ZN(new_n753));
  AOI211_X1 g552(.A(KEYINPUT87), .B(new_n579), .C1(new_n581), .C2(new_n585), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n748), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n589), .A2(KEYINPUT100), .A3(new_n746), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(KEYINPUT101), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n752), .A2(new_n758), .A3(new_n744), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(KEYINPUT102), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT102), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n750), .B1(new_n761), .B2(new_n762), .ZN(G1330gat));
  NAND3_X1  g562(.A1(new_n724), .A2(new_n387), .A3(new_n725), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(new_n767), .A3(new_n515), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n730), .A2(new_n515), .A3(new_n387), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(KEYINPUT48), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(G50gat), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n769), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT103), .B(KEYINPUT48), .Z(new_n775));
  OAI22_X1  g574(.A1(new_n768), .A2(new_n772), .B1(new_n774), .B2(new_n775), .ZN(G1331gat));
  INV_X1    g575(.A(new_n663), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n579), .A2(new_n686), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n508), .A2(new_n777), .A3(new_n718), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n695), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(new_n641), .Z(G1332gat));
  AOI21_X1  g580(.A(new_n465), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT106), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT107), .Z(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1333gat));
  NAND2_X1  g586(.A1(new_n779), .A2(new_n742), .ZN(new_n788));
  INV_X1    g587(.A(new_n501), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(G71gat), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n788), .A2(G71gat), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1334gat));
  NAND2_X1  g592(.A1(new_n779), .A2(new_n387), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g594(.A1(new_n578), .A2(new_n663), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT109), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n686), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n724), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n439), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n720), .A2(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n803), .A2(new_n592), .A3(new_n695), .A4(new_n686), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n687), .A2(new_n465), .A3(G92gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n798), .A2(new_n721), .A3(new_n464), .A4(new_n723), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n802), .A2(KEYINPUT111), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n815), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n811), .B1(new_n818), .B2(new_n813), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n808), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n818), .A2(new_n813), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(KEYINPUT112), .C1(new_n822), .C2(new_n811), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n799), .B2(new_n705), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n789), .A2(G99gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n803), .A2(new_n686), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1338gat));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g628(.A(G106gat), .B1(new_n799), .B2(new_n503), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n687), .A2(new_n503), .A3(G106gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n803), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n829), .B(new_n830), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n816), .B2(new_n817), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT53), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(G1339gat));
  NAND3_X1  g638(.A1(new_n667), .A2(new_n674), .A3(new_n666), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n680), .B1(new_n675), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n685), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(new_n841), .B2(new_n843), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n576), .B2(new_n577), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n556), .A2(new_n561), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n573), .A2(new_n548), .B1(new_n850), .B2(new_n560), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n570), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n575), .A2(new_n686), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n635), .A3(new_n664), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n848), .A2(new_n575), .A3(new_n852), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n627), .A2(new_n633), .A3(new_n631), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n633), .B1(new_n627), .B2(new_n631), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n663), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n688), .A2(new_n578), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n506), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n439), .A2(new_n464), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n579), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(new_n259), .ZN(G1340gat));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n687), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(new_n257), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n663), .A3(new_n864), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n252), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n252), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n873), .B2(new_n872), .ZN(G1342gat));
  NAND2_X1  g674(.A1(new_n855), .A2(new_n859), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n777), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n689), .A2(new_n579), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n506), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n718), .A4(new_n864), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n881), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT115), .B1(new_n881), .B2(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(G134gat), .B1(new_n881), .B2(KEYINPUT56), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n884), .B(new_n885), .Z(G1343gat));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  INV_X1    g686(.A(new_n864), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n742), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n862), .B2(new_n503), .ZN(new_n892));
  INV_X1    g691(.A(new_n853), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n894));
  XNOR2_X1  g693(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n844), .B2(KEYINPUT116), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n846), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n893), .B1(new_n578), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n859), .B1(new_n718), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n777), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n878), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n503), .A2(new_n891), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n890), .B1(new_n892), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n579), .A2(new_n332), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n879), .A2(new_n387), .A3(new_n889), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(G141gat), .B1(new_n908), .B2(new_n578), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n887), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n887), .B(new_n912), .C1(new_n906), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n333), .A3(new_n686), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n387), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n891), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n879), .A2(new_n902), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n686), .A3(new_n889), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n916), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT59), .B(new_n333), .C1(new_n904), .C2(new_n686), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(G1345gat));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n329), .A3(new_n663), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n904), .A2(new_n663), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n329), .ZN(G1346gat));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n320), .A3(new_n718), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n904), .A2(new_n718), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n320), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n695), .A2(new_n465), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n880), .B(new_n931), .C1(new_n860), .C2(new_n861), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n203), .A3(new_n578), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n879), .A2(KEYINPUT119), .A3(new_n880), .A4(new_n931), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n578), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT120), .A3(G169gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT120), .B1(new_n939), .B2(G169gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(G1348gat));
  OAI21_X1  g741(.A(new_n204), .B1(new_n932), .B2(new_n687), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT121), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n687), .A2(new_n204), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n938), .B2(new_n945), .ZN(G1349gat));
  NAND2_X1  g745(.A1(new_n663), .A2(new_n212), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n932), .A2(new_n947), .B1(KEYINPUT123), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(KEYINPUT123), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n937), .A3(new_n663), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n238), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT122), .A4(new_n663), .ZN(new_n955));
  AOI211_X1 g754(.A(new_n949), .B(new_n951), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n952), .A2(new_n953), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(G183gat), .A3(new_n955), .ZN(new_n958));
  INV_X1    g757(.A(new_n949), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n956), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n933), .A2(new_n213), .A3(new_n718), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n938), .A2(new_n718), .ZN(new_n963));
  XNOR2_X1  g762(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n963), .A2(G190gat), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n963), .B2(G190gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  NAND2_X1  g766(.A1(new_n931), .A2(new_n387), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n862), .A2(new_n742), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(G197gat), .B1(new_n969), .B2(new_n578), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n705), .A2(new_n931), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n918), .B2(new_n919), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n578), .A2(G197gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  INV_X1    g773(.A(G204gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n972), .B2(new_n686), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n742), .A2(new_n968), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n879), .A2(new_n975), .A3(new_n686), .A4(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n981), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(KEYINPUT126), .B1(new_n976), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n981), .B(new_n982), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  AOI211_X1 g786(.A(new_n687), .B(new_n971), .C1(new_n918), .C2(new_n919), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n986), .B(new_n987), .C1(new_n975), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n985), .A2(new_n989), .ZN(G1353gat));
  INV_X1    g789(.A(G211gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n969), .A2(new_n991), .A3(new_n663), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n972), .A2(new_n663), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995));
  AOI211_X1 g794(.A(new_n995), .B(new_n991), .C1(new_n972), .C2(new_n663), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n994), .B2(new_n996), .ZN(G1354gat));
  AOI21_X1  g796(.A(G218gat), .B1(new_n969), .B2(new_n718), .ZN(new_n998));
  OR2_X1    g797(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n719), .A2(new_n590), .ZN(new_n1001));
  AOI22_X1  g800(.A1(new_n999), .A2(new_n1000), .B1(new_n972), .B2(new_n1001), .ZN(G1355gat));
endmodule


