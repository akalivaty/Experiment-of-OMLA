//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT64), .A3(G143), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G146), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n195), .A2(new_n197), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G104), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(G107), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n196), .A2(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n198), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT68), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n200), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n201), .B(new_n213), .C1(new_n217), .C2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n195), .A2(new_n197), .A3(new_n200), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n201), .B1(new_n224), .B2(new_n215), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n209), .A2(new_n212), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G134), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(G134), .A3(new_n230), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n230), .A2(G134), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G137), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n237), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n244), .A3(new_n234), .A4(new_n233), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n233), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n228), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n228), .B(new_n249), .C1(new_n251), .C2(KEYINPUT12), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n203), .A2(new_n206), .A3(new_n208), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT76), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n203), .A2(new_n206), .A3(new_n259), .A4(new_n208), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  OR2_X1    g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n221), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n195), .A2(new_n197), .A3(new_n266), .A4(new_n200), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n258), .A2(G101), .A3(new_n260), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT10), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n269), .A2(new_n271), .B1(new_n272), .B2(new_n227), .ZN(new_n273));
  INV_X1    g087(.A(new_n201), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT68), .B1(new_n215), .B2(new_n216), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n220), .A2(new_n218), .A3(new_n221), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n209), .A2(new_n212), .A3(KEYINPUT10), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT77), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n201), .B1(new_n217), .B2(new_n222), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n281));
  INV_X1    g095(.A(new_n278), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n240), .A2(new_n245), .B1(G131), .B2(new_n247), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n273), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n192), .B1(new_n256), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n273), .B2(new_n284), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n286), .A2(new_n192), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n187), .B(G469), .C1(new_n291), .C2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(G469), .A2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n273), .A2(new_n284), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n295), .A2(new_n285), .B1(new_n254), .B2(new_n255), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n286), .A2(new_n192), .ZN(new_n297));
  OAI22_X1  g111(.A1(new_n296), .A2(new_n192), .B1(new_n288), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT79), .B(new_n293), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(KEYINPUT80), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n286), .A2(new_n303), .A3(new_n192), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n304), .A3(new_n256), .ZN(new_n305));
  INV_X1    g119(.A(new_n286), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n191), .B1(new_n306), .B2(new_n288), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n299), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n299), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT81), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n301), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(G116), .B(G119), .Z(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n271), .A2(new_n318), .A3(new_n262), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G116), .ZN(new_n323));
  OAI211_X1 g137(.A(G113), .B(new_n323), .C1(new_n316), .C2(new_n321), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n226), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(G110), .B(G122), .Z(new_n327));
  OR2_X1    g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT6), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n277), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n265), .A2(new_n267), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n189), .A2(G224), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n335), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n326), .A2(new_n339), .A3(new_n327), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n330), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n324), .A2(new_n320), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n213), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n325), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n327), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n335), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(new_n336), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT7), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n335), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT7), .B1(new_n336), .B2(KEYINPUT83), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(KEYINPUT83), .B2(new_n336), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n332), .A2(new_n334), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT84), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n337), .A2(new_n335), .B1(new_n344), .B2(new_n346), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT84), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n351), .A4(new_n354), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n359), .A3(new_n328), .ZN(new_n360));
  INV_X1    g174(.A(G902), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n341), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G210), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n341), .A2(new_n360), .A3(new_n361), .A4(new_n363), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n315), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(G221), .B1(new_n369), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G125), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n331), .A2(G140), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT73), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(KEYINPUT73), .A3(G125), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G146), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n196), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n379), .B1(new_n378), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  AND4_X1   g199(.A1(G143), .A2(new_n385), .A3(new_n189), .A4(G214), .ZN(new_n386));
  NOR2_X1   g200(.A1(G237), .A2(G953), .ZN(new_n387));
  AOI21_X1  g201(.A(G143), .B1(new_n387), .B2(G214), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT18), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(KEYINPUT86), .C1(new_n390), .C2(new_n234), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n189), .A3(G214), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n194), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n393), .B(new_n394), .C1(new_n390), .C2(new_n234), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n234), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT18), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n384), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n202), .ZN(new_n403));
  INV_X1    g217(.A(new_n398), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n389), .A2(new_n234), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n377), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n373), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G146), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n196), .A3(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n398), .A2(KEYINPUT17), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n407), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n401), .A2(new_n403), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n403), .B1(new_n401), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n361), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G475), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n380), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n376), .A2(new_n377), .B1(new_n380), .B2(KEYINPUT87), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n196), .B(new_n424), .C1(new_n425), .C2(new_n423), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n412), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT88), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n412), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n404), .A2(new_n405), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n403), .B1(new_n432), .B2(new_n401), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n420), .B(new_n421), .C1(new_n433), .C2(new_n416), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n401), .A2(new_n403), .A3(new_n415), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n384), .A2(new_n400), .ZN(new_n437));
  INV_X1    g251(.A(new_n431), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n427), .B2(KEYINPUT88), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n440), .B2(new_n403), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n420), .B1(new_n441), .B2(new_n421), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n419), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT89), .B(new_n419), .C1(new_n435), .C2(new_n442), .ZN(new_n446));
  INV_X1    g260(.A(G234), .ZN(new_n447));
  OAI211_X1 g261(.A(G952), .B(new_n189), .C1(new_n447), .C2(new_n385), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n448), .B(KEYINPUT92), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(G902), .B(G953), .C1(new_n447), .C2(new_n385), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT93), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G478), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT13), .B1(new_n198), .B2(G143), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n241), .ZN(new_n461));
  XNOR2_X1  g275(.A(G128), .B(G143), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G116), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT90), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(G107), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(G107), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n469));
  INV_X1    g283(.A(G116), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(G122), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT91), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n205), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT91), .B1(new_n472), .B2(KEYINPUT14), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n462), .B(new_n241), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n478), .C1(G107), .C2(new_n465), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n369), .A2(new_n481), .A3(G953), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n480), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n459), .B1(new_n484), .B2(new_n361), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n483), .A2(G902), .A3(new_n458), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n445), .A2(new_n446), .A3(new_n456), .A4(new_n487), .ZN(new_n488));
  NOR4_X1   g302(.A1(new_n313), .A2(new_n368), .A3(new_n371), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n412), .ZN(new_n490));
  INV_X1    g304(.A(new_n381), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n322), .B2(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n322), .A2(G128), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G110), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT24), .B(G110), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n322), .A2(KEYINPUT72), .A3(G128), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT72), .B1(new_n322), .B2(G128), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n494), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OR3_X1    g316(.A1(new_n490), .A2(new_n491), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(G110), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n501), .B2(new_n498), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n412), .B2(new_n413), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT22), .B(G137), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n510), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n490), .A2(new_n502), .A3(new_n491), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n506), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n481), .B1(G234), .B2(new_n361), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n361), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT75), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n514), .A3(new_n361), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT25), .A4(new_n361), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n517), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G472), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n242), .B2(new_n237), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT67), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n246), .A2(new_n280), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n333), .B1(new_n246), .B2(new_n248), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n318), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n246), .A2(new_n280), .A3(new_n532), .ZN(new_n536));
  INV_X1    g350(.A(new_n318), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(new_n285), .C2(new_n333), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n530), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n530), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n387), .A2(G210), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT29), .ZN(new_n547));
  INV_X1    g361(.A(new_n538), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n533), .B2(new_n534), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n536), .B(KEYINPUT30), .C1(new_n285), .C2(new_n333), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n318), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT69), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n550), .A2(KEYINPUT69), .A3(new_n318), .A4(new_n551), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n547), .B1(new_n556), .B2(new_n544), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n546), .B2(KEYINPUT29), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n529), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n538), .A2(new_n544), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n554), .B2(new_n555), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n545), .B1(new_n539), .B2(new_n540), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT71), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n572), .B(new_n545), .C1(new_n539), .C2(new_n540), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n564), .A2(new_n568), .A3(new_n569), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n559), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n528), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n489), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  NOR3_X1   g397(.A1(new_n313), .A2(new_n528), .A3(new_n371), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n367), .A2(new_n456), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n445), .A2(new_n446), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n484), .A2(KEYINPUT33), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n483), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(G478), .B(new_n361), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT94), .B(G478), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n483), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n577), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n529), .B1(new_n575), .B2(new_n361), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  INV_X1    g416(.A(new_n487), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n435), .A2(new_n442), .A3(KEYINPUT95), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n442), .A2(KEYINPUT95), .B1(G475), .B2(new_n418), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n602), .B1(new_n585), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n608), .A2(new_n367), .A3(KEYINPUT96), .A4(new_n456), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n584), .A3(new_n598), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n503), .A2(new_n507), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n519), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n614), .B1(new_n619), .B2(new_n526), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n527), .A2(KEYINPUT97), .A3(new_n618), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n367), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n596), .A2(new_n622), .A3(new_n597), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n313), .A2(new_n371), .A3(new_n488), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  NAND2_X1  g441(.A1(new_n577), .A2(new_n578), .ZN(new_n628));
  INV_X1    g442(.A(new_n559), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n580), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n313), .A2(new_n371), .ZN(new_n631));
  INV_X1    g445(.A(new_n622), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n450), .B1(new_n633), .B2(new_n453), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n606), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n630), .A2(new_n631), .A3(new_n632), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  XOR2_X1   g451(.A(new_n634), .B(KEYINPUT39), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT40), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n365), .A2(new_n366), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n641), .B(new_n642), .Z(new_n643));
  NAND2_X1  g457(.A1(new_n586), .A2(new_n603), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n643), .A2(new_n315), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n619), .A2(new_n526), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n544), .B1(new_n535), .B2(new_n538), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n563), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n529), .B1(new_n650), .B2(new_n361), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n577), .B2(new_n578), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n647), .B1(new_n652), .B2(new_n580), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n640), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n194), .ZN(G45));
  NOR2_X1   g470(.A1(new_n594), .A2(new_n634), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n630), .A2(new_n631), .A3(new_n632), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NAND2_X1  g473(.A1(new_n312), .A2(new_n310), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n299), .B1(new_n308), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n661), .B2(new_n308), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n371), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n581), .A2(new_n595), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND3_X1  g482(.A1(new_n581), .A2(new_n610), .A3(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  INV_X1    g484(.A(new_n586), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n621), .A2(new_n620), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n603), .A2(new_n455), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n579), .B2(new_n580), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n660), .A2(new_n663), .A3(new_n370), .A4(new_n367), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  INV_X1    g493(.A(new_n528), .ZN(new_n680));
  INV_X1    g494(.A(new_n576), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n539), .A2(new_n540), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n563), .A2(KEYINPUT31), .B1(new_n545), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n681), .B1(new_n683), .B2(new_n569), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n575), .A2(new_n361), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n680), .B(new_n685), .C1(new_n686), .C2(new_n529), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n586), .B2(new_n603), .ZN(new_n689));
  AOI211_X1 g503(.A(KEYINPUT101), .B(new_n487), .C1(new_n445), .C2(new_n446), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n676), .A2(new_n455), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  NOR3_X1   g509(.A1(new_n597), .A2(new_n646), .A3(new_n684), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n677), .A2(new_n696), .A3(new_n657), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n575), .A2(KEYINPUT105), .A3(KEYINPUT32), .A4(new_n576), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n580), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n579), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n680), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n305), .A2(new_n307), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n309), .A2(new_n705), .A3(new_n299), .A4(new_n361), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n309), .B1(new_n308), .B2(new_n299), .ZN(new_n707));
  AOI211_X1 g521(.A(KEYINPUT102), .B(new_n192), .C1(new_n256), .C2(new_n286), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n253), .B1(new_n285), .B2(KEYINPUT78), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n227), .A2(new_n223), .B1(new_n246), .B2(new_n248), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n255), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n286), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n709), .B1(new_n714), .B2(new_n191), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n290), .A2(KEYINPUT103), .A3(new_n289), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n297), .B2(new_n288), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(G902), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  OAI22_X1  g535(.A1(new_n706), .A2(new_n707), .B1(new_n721), .B2(new_n299), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT102), .B1(new_n296), .B2(new_n192), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n287), .A2(new_n709), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n720), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n361), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(KEYINPUT104), .C1(new_n706), .C2(new_n707), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n370), .A2(new_n314), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n641), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n634), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n586), .A2(KEYINPUT42), .A3(new_n593), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n731), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n699), .B1(new_n704), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g553(.A(new_n733), .B(new_n736), .C1(new_n724), .C2(new_n730), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n680), .A4(new_n703), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n733), .B1(new_n724), .B2(new_n730), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n581), .A2(new_n743), .A3(new_n657), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n739), .A2(new_n741), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n234), .ZN(G33));
  NAND3_X1  g560(.A1(new_n581), .A2(new_n743), .A3(new_n635), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n586), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n593), .A2(KEYINPUT43), .ZN(new_n751));
  INV_X1    g565(.A(new_n593), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n586), .ZN(new_n753));
  OAI22_X1  g567(.A1(new_n750), .A2(new_n751), .B1(KEYINPUT43), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n598), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n647), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT108), .Z(new_n759));
  NAND3_X1  g573(.A1(new_n365), .A2(new_n314), .A3(new_n366), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n716), .A2(KEYINPUT45), .A3(new_n720), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(G469), .C1(KEYINPUT45), .C2(new_n291), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n293), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n660), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n370), .A3(new_n638), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n760), .B(new_n769), .C1(new_n756), .C2(new_n757), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n759), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(G137), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G39));
  INV_X1    g587(.A(new_n760), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n657), .A2(new_n528), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n630), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT47), .B1(new_n768), .B2(new_n370), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT47), .B(new_n370), .C1(new_n766), .C2(new_n767), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n776), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  INV_X1    g595(.A(new_n643), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n782), .A2(new_n528), .A3(new_n752), .A4(new_n732), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n652), .A2(new_n580), .ZN(new_n784));
  INV_X1    g598(.A(new_n750), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n664), .B(KEYINPUT49), .Z(new_n786));
  NAND4_X1  g600(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n636), .A2(new_n658), .A3(new_n697), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n735), .A2(KEYINPUT113), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n735), .A2(KEYINPUT113), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n791), .A3(new_n371), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n724), .B2(new_n730), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n644), .A2(KEYINPUT101), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n586), .A2(new_n688), .A3(new_n603), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n368), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n653), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n789), .A2(new_n799), .A3(KEYINPUT114), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n636), .A2(new_n658), .A3(new_n697), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n798), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n789), .B2(new_n799), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n672), .A2(new_n487), .A3(new_n735), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n604), .A2(new_n605), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(new_n760), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n630), .A3(new_n631), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n743), .A2(new_n657), .A3(new_n696), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n747), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT111), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n747), .A2(new_n812), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n692), .A2(new_n693), .B1(new_n675), .B2(new_n677), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n489), .A2(new_n581), .B1(new_n623), .B2(new_n624), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n671), .A2(KEYINPUT110), .A3(new_n603), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n586), .B2(new_n487), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n594), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n585), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n584), .A3(new_n825), .A4(new_n598), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n581), .B(new_n665), .C1(new_n610), .C2(new_n595), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n819), .A2(new_n820), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n739), .A2(new_n741), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n744), .A2(new_n742), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n808), .A2(new_n818), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n745), .A2(new_n828), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n808), .B1(new_n834), .B2(new_n818), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n788), .B(new_n807), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT114), .B1(new_n789), .B2(new_n799), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n802), .A2(new_n798), .A3(new_n801), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n805), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n800), .A2(KEYINPUT52), .A3(new_n803), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n818), .A2(new_n829), .A3(new_n832), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT112), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n834), .A2(new_n808), .A3(new_n818), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n836), .B(KEYINPUT54), .C1(new_n845), .C2(new_n788), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n807), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n834), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n848), .B(new_n849), .C1(new_n845), .C2(KEYINPUT53), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n846), .B2(new_n850), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  INV_X1    g667(.A(new_n664), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n733), .A2(new_n449), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n754), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n680), .A2(new_n784), .A3(new_n854), .A4(new_n855), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n586), .A2(new_n593), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n856), .A2(new_n696), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n664), .A2(new_n370), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n777), .A2(new_n779), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n687), .A2(new_n449), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n754), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(new_n774), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(KEYINPUT116), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(KEYINPUT116), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n665), .A2(new_n315), .A3(new_n643), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT50), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n863), .A2(KEYINPUT50), .A3(new_n869), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n853), .B1(new_n868), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n704), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n856), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n863), .A2(new_n677), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n189), .A2(G952), .ZN(new_n885));
  INV_X1    g699(.A(new_n594), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n857), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n865), .A2(KEYINPUT51), .A3(new_n859), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n882), .B(new_n888), .C1(new_n889), .C2(new_n876), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n878), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n851), .A2(new_n852), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n787), .B1(new_n892), .B2(new_n893), .ZN(G75));
  OAI21_X1  g708(.A(new_n849), .B1(new_n845), .B2(KEYINPUT53), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(G210), .A3(G902), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n330), .A2(new_n340), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n338), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n896), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n896), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n189), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  XOR2_X1   g719(.A(new_n293), .B(KEYINPUT57), .Z(new_n906));
  INV_X1    g720(.A(new_n840), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n804), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n833), .B2(new_n835), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n788), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n848), .B1(new_n910), .B2(new_n849), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n818), .A2(new_n829), .A3(new_n832), .A4(KEYINPUT53), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n804), .A3(new_n806), .ZN(new_n913));
  AOI211_X1 g727(.A(KEYINPUT54), .B(new_n913), .C1(new_n909), .C2(new_n788), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n705), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n762), .B(KEYINPUT121), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n895), .A2(G902), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n904), .B1(new_n916), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n843), .A2(new_n844), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n921), .B2(new_n908), .ZN(new_n922));
  OAI211_X1 g736(.A(G902), .B(new_n920), .C1(new_n922), .C2(new_n913), .ZN(new_n923));
  INV_X1    g737(.A(new_n441), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n904), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n895), .A2(G902), .A3(new_n441), .A4(new_n920), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n926), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(G60));
  OR2_X1    g746(.A1(new_n587), .A2(new_n589), .ZN(new_n933));
  XOR2_X1   g747(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n457), .A2(new_n361), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n911), .B2(new_n914), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n926), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n851), .B2(new_n852), .ZN(new_n940));
  INV_X1    g754(.A(new_n933), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n910), .B2(new_n849), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(new_n515), .ZN(new_n946));
  INV_X1    g760(.A(new_n944), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n895), .A2(new_n617), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n926), .A4(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(new_n926), .C1(new_n945), .C2(new_n515), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(G66));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n454), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n829), .B2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n897), .B1(G898), .B2(new_n189), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  NOR2_X1   g772(.A1(new_n655), .A2(new_n802), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  INV_X1    g774(.A(new_n639), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n581), .A3(new_n774), .A4(new_n824), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n780), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n759), .B2(new_n770), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n189), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n550), .A2(new_n551), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n424), .B1(new_n425), .B2(new_n423), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  AOI21_X1  g786(.A(G953), .B1(new_n960), .B2(new_n964), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n969), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n769), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n879), .A3(new_n797), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n747), .A2(new_n980), .A3(new_n780), .A4(new_n789), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n771), .A2(new_n981), .A3(new_n832), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n189), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n983), .A2(new_n984), .B1(new_n977), .B2(new_n976), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n975), .A2(new_n978), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n978), .B1(new_n975), .B2(new_n985), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G72));
  NOR2_X1   g803(.A1(new_n556), .A2(new_n545), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n965), .A2(new_n828), .ZN(new_n991));
  XNOR2_X1  g805(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n529), .A2(new_n361), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n992), .B(new_n993), .Z(new_n994));
  OAI21_X1  g808(.A(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n556), .A2(new_n545), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n982), .B2(new_n829), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n995), .B(new_n926), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n836), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(KEYINPUT53), .B2(new_n909), .ZN(new_n1000));
  INV_X1    g814(.A(new_n996), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n1001), .A2(new_n990), .A3(new_n994), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT127), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1000), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n998), .B1(new_n1004), .B2(new_n1006), .ZN(G57));
endmodule


