

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797;

  XNOR2_X1 U371 ( .A(n403), .B(KEYINPUT105), .ZN(n402) );
  XNOR2_X1 U372 ( .A(n518), .B(n517), .ZN(n774) );
  XNOR2_X1 U373 ( .A(G116), .B(G119), .ZN(n471) );
  NAND2_X2 U374 ( .A1(n492), .A2(n680), .ZN(n695) );
  NAND2_X2 U375 ( .A1(n421), .A2(KEYINPUT1), .ZN(n406) );
  OR2_X2 U376 ( .A1(n567), .A2(n586), .ZN(n569) );
  XNOR2_X2 U377 ( .A(n593), .B(KEYINPUT104), .ZN(n612) );
  XNOR2_X2 U378 ( .A(n392), .B(KEYINPUT40), .ZN(n633) );
  BUF_X2 U379 ( .A(n594), .Z(n596) );
  XNOR2_X2 U380 ( .A(n774), .B(n528), .ZN(n685) );
  XNOR2_X2 U381 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n368) );
  XNOR2_X2 U382 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X2 U383 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X2 U384 ( .A(n593), .B(n419), .ZN(n607) );
  NOR2_X2 U385 ( .A1(n653), .A2(n652), .ZN(n452) );
  INV_X1 U386 ( .A(n492), .ZN(n479) );
  XOR2_X1 U387 ( .A(n543), .B(n542), .Z(n350) );
  AND2_X2 U388 ( .A1(n461), .A2(n456), .ZN(n455) );
  NOR2_X2 U389 ( .A1(n724), .A2(n726), .ZN(n747) );
  INV_X2 U390 ( .A(n731), .ZN(n351) );
  XNOR2_X2 U391 ( .A(G953), .B(KEYINPUT64), .ZN(n492) );
  NAND2_X1 U392 ( .A1(n660), .A2(n724), .ZN(n392) );
  XNOR2_X1 U393 ( .A(n423), .B(n628), .ZN(n660) );
  AND2_X1 U394 ( .A1(n638), .A2(n637), .ZN(n641) );
  AND2_X1 U395 ( .A1(n624), .A2(n626), .ZN(n433) );
  NAND2_X2 U396 ( .A1(n430), .A2(n386), .ZN(n421) );
  BUF_X1 U397 ( .A(n706), .Z(n352) );
  INV_X1 U398 ( .A(n664), .ZN(n353) );
  BUF_X1 U399 ( .A(n618), .Z(n592) );
  NOR2_X2 U400 ( .A1(n648), .A2(n753), .ZN(n533) );
  BUF_X1 U401 ( .A(n537), .Z(n354) );
  NOR2_X1 U402 ( .A1(n618), .A2(KEYINPUT44), .ZN(n439) );
  XNOR2_X2 U403 ( .A(n537), .B(KEYINPUT4), .ZN(n525) );
  XNOR2_X2 U404 ( .A(n467), .B(G128), .ZN(n537) );
  XNOR2_X2 U405 ( .A(n503), .B(n366), .ZN(n417) );
  NOR2_X1 U406 ( .A1(n376), .A2(n378), .ZN(n639) );
  NAND2_X1 U407 ( .A1(n355), .A2(n379), .ZN(n378) );
  XNOR2_X1 U408 ( .A(n523), .B(n411), .ZN(n547) );
  XNOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n411) );
  XNOR2_X1 U410 ( .A(n559), .B(n558), .ZN(n591) );
  XOR2_X1 U411 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n549) );
  INV_X1 U412 ( .A(KEYINPUT108), .ZN(n385) );
  XNOR2_X1 U413 ( .A(n409), .B(n486), .ZN(n487) );
  NOR2_X1 U414 ( .A1(G953), .A2(G237), .ZN(n550) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n468) );
  INV_X1 U416 ( .A(KEYINPUT34), .ZN(n448) );
  AND2_X1 U417 ( .A1(n351), .A2(n385), .ZN(n381) );
  NOR2_X1 U418 ( .A1(n384), .A2(n383), .ZN(n382) );
  NOR2_X1 U419 ( .A1(n351), .A2(n385), .ZN(n384) );
  NOR2_X1 U420 ( .A1(n514), .A2(n385), .ZN(n383) );
  INV_X1 U421 ( .A(KEYINPUT3), .ZN(n470) );
  XNOR2_X1 U422 ( .A(G128), .B(G110), .ZN(n482) );
  NAND2_X1 U423 ( .A1(n397), .A2(n395), .ZN(n535) );
  AND2_X1 U424 ( .A1(n400), .A2(n398), .ZN(n397) );
  NAND2_X1 U425 ( .A1(n479), .A2(n396), .ZN(n395) );
  NAND2_X1 U426 ( .A1(n480), .A2(n399), .ZN(n398) );
  XNOR2_X1 U427 ( .A(n547), .B(n485), .ZN(n785) );
  XNOR2_X1 U428 ( .A(n422), .B(n557), .ZN(n692) );
  XNOR2_X1 U429 ( .A(n547), .B(n358), .ZN(n422) );
  XNOR2_X1 U430 ( .A(G107), .B(KEYINPUT78), .ZN(n508) );
  XOR2_X1 U431 ( .A(G104), .B(G110), .Z(n509) );
  NAND2_X1 U432 ( .A1(n433), .A2(n434), .ZN(n423) );
  INV_X1 U433 ( .A(KEYINPUT6), .ZN(n419) );
  XNOR2_X1 U434 ( .A(n580), .B(n579), .ZN(n610) );
  XNOR2_X1 U435 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n579) );
  NOR2_X1 U436 ( .A1(n729), .A2(n544), .ZN(n442) );
  NAND2_X1 U437 ( .A1(G469), .A2(n429), .ZN(n428) );
  NAND2_X1 U438 ( .A1(n513), .A2(G902), .ZN(n431) );
  XNOR2_X1 U439 ( .A(n410), .B(KEYINPUT20), .ZN(n497) );
  INV_X1 U440 ( .A(G234), .ZN(n399) );
  INV_X1 U441 ( .A(KEYINPUT8), .ZN(n480) );
  NOR2_X1 U442 ( .A1(n480), .A2(n399), .ZN(n396) );
  INV_X1 U443 ( .A(KEYINPUT65), .ZN(n462) );
  NAND2_X1 U444 ( .A1(n458), .A2(n457), .ZN(n456) );
  NAND2_X1 U445 ( .A1(n460), .A2(n459), .ZN(n458) );
  NAND2_X1 U446 ( .A1(KEYINPUT2), .A2(KEYINPUT65), .ZN(n459) );
  XNOR2_X1 U447 ( .A(G122), .B(G113), .ZN(n548) );
  XNOR2_X1 U448 ( .A(G143), .B(G104), .ZN(n553) );
  XOR2_X1 U449 ( .A(G140), .B(G131), .Z(n554) );
  INV_X1 U450 ( .A(KEYINPUT92), .ZN(n519) );
  XOR2_X1 U451 ( .A(G146), .B(G125), .Z(n523) );
  NAND2_X1 U452 ( .A1(G237), .A2(G234), .ZN(n490) );
  OR2_X1 U453 ( .A1(G902), .A2(G237), .ZN(n531) );
  XNOR2_X1 U454 ( .A(G107), .B(G134), .ZN(n538) );
  XOR2_X1 U455 ( .A(G122), .B(G116), .Z(n539) );
  AND2_X1 U456 ( .A1(n563), .A2(n664), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n435), .B(n368), .ZN(n618) );
  INV_X1 U458 ( .A(n647), .ZN(n447) );
  XNOR2_X1 U459 ( .A(n373), .B(n372), .ZN(n741) );
  INV_X1 U460 ( .A(KEYINPUT98), .ZN(n372) );
  XNOR2_X1 U461 ( .A(n375), .B(KEYINPUT77), .ZN(n374) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n624) );
  INV_X1 U463 ( .A(KEYINPUT30), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n622), .B(KEYINPUT79), .ZN(n434) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n600) );
  XNOR2_X1 U466 ( .A(n544), .B(KEYINPUT103), .ZN(n404) );
  NAND2_X1 U467 ( .A1(n350), .A2(n429), .ZN(n405) );
  INV_X1 U468 ( .A(n788), .ZN(n418) );
  INV_X1 U469 ( .A(KEYINPUT16), .ZN(n425) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n412) );
  NAND2_X1 U471 ( .A1(n535), .A2(G221), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n484), .B(n481), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n415), .B(n370), .ZN(n795) );
  NOR2_X1 U474 ( .A1(n610), .A2(n609), .ZN(n415) );
  AND2_X1 U475 ( .A1(n599), .A2(n600), .ZN(n726) );
  XNOR2_X1 U476 ( .A(n446), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U477 ( .A(n443), .B(n350), .ZN(n424) );
  NAND2_X1 U478 ( .A1(n442), .A2(n441), .ZN(n443) );
  XNOR2_X1 U479 ( .A(n633), .B(G131), .ZN(G33) );
  AND2_X1 U480 ( .A1(n416), .A2(n514), .ZN(n355) );
  INV_X1 U481 ( .A(G902), .ZN(n429) );
  NOR2_X1 U482 ( .A1(n734), .A2(n500), .ZN(n356) );
  AND2_X1 U483 ( .A1(n643), .A2(n642), .ZN(n357) );
  XOR2_X1 U484 ( .A(n546), .B(n545), .Z(n358) );
  INV_X1 U485 ( .A(n747), .ZN(n379) );
  AND2_X1 U486 ( .A1(n427), .A2(n463), .ZN(n359) );
  NOR2_X1 U487 ( .A1(n636), .A2(n747), .ZN(n360) );
  AND2_X1 U488 ( .A1(n514), .A2(n351), .ZN(n361) );
  AND2_X1 U489 ( .A1(n382), .A2(n380), .ZN(n362) );
  AND2_X1 U490 ( .A1(n357), .A2(n355), .ZN(n363) );
  AND2_X1 U491 ( .A1(n363), .A2(n417), .ZN(n364) );
  AND2_X1 U492 ( .A1(n402), .A2(n563), .ZN(n365) );
  XOR2_X1 U493 ( .A(n502), .B(n501), .Z(n366) );
  XOR2_X1 U494 ( .A(KEYINPUT66), .B(KEYINPUT19), .Z(n367) );
  OR2_X1 U495 ( .A1(n671), .A2(n462), .ZN(n369) );
  XOR2_X1 U496 ( .A(KEYINPUT80), .B(KEYINPUT32), .Z(n370) );
  XNOR2_X1 U497 ( .A(n412), .B(n785), .ZN(n700) );
  INV_X1 U498 ( .A(KEYINPUT2), .ZN(n463) );
  AND2_X1 U499 ( .A1(n463), .A2(n462), .ZN(n371) );
  NAND2_X1 U500 ( .A1(n374), .A2(n593), .ZN(n373) );
  NAND2_X1 U501 ( .A1(n407), .A2(n406), .ZN(n375) );
  INV_X1 U502 ( .A(n417), .ZN(n376) );
  INV_X1 U503 ( .A(n377), .ZN(n534) );
  NAND2_X1 U504 ( .A1(n417), .A2(n355), .ZN(n377) );
  NAND2_X1 U505 ( .A1(n381), .A2(n514), .ZN(n380) );
  XNOR2_X2 U506 ( .A(n595), .B(KEYINPUT31), .ZN(n727) );
  NAND2_X1 U507 ( .A1(n736), .A2(n420), .ZN(n737) );
  NAND2_X1 U508 ( .A1(n361), .A2(n420), .ZN(n597) );
  NAND2_X1 U509 ( .A1(n607), .A2(n356), .ZN(n403) );
  XNOR2_X1 U510 ( .A(n533), .B(n367), .ZN(n416) );
  XNOR2_X1 U511 ( .A(n473), .B(n472), .ZN(n515) );
  XNOR2_X1 U512 ( .A(n515), .B(n425), .ZN(n518) );
  OR2_X1 U513 ( .A1(n706), .A2(n428), .ZN(n386) );
  NOR2_X1 U514 ( .A1(n388), .A2(KEYINPUT1), .ZN(n387) );
  NOR2_X1 U515 ( .A1(n706), .A2(n428), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n407), .A2(n406), .ZN(n389) );
  BUF_X1 U517 ( .A(n408), .Z(n390) );
  INV_X1 U518 ( .A(n421), .ZN(n514) );
  NAND2_X1 U519 ( .A1(n497), .A2(G217), .ZN(n409) );
  XNOR2_X1 U520 ( .A(n489), .B(n488), .ZN(n585) );
  BUF_X1 U521 ( .A(n585), .Z(n734) );
  XNOR2_X1 U522 ( .A(n389), .B(KEYINPUT77), .ZN(n453) );
  NAND2_X1 U523 ( .A1(n745), .A2(n594), .ZN(n590) );
  XNOR2_X1 U524 ( .A(n589), .B(n588), .ZN(n745) );
  NAND2_X1 U525 ( .A1(n612), .A2(n356), .ZN(n503) );
  NAND2_X1 U526 ( .A1(n612), .A2(n623), .ZN(n394) );
  XOR2_X1 U527 ( .A(KEYINPUT62), .B(n677), .Z(n678) );
  NAND2_X1 U528 ( .A1(n455), .A2(n454), .ZN(n676) );
  INV_X1 U529 ( .A(n676), .ZN(n441) );
  XNOR2_X1 U530 ( .A(n391), .B(n659), .ZN(n670) );
  NAND2_X1 U531 ( .A1(n657), .A2(n658), .ZN(n391) );
  NOR2_X2 U532 ( .A1(n727), .A2(n713), .ZN(n601) );
  NAND2_X1 U533 ( .A1(n492), .A2(n480), .ZN(n400) );
  NAND2_X1 U534 ( .A1(n401), .A2(n402), .ZN(n566) );
  NAND2_X1 U535 ( .A1(n387), .A2(n430), .ZN(n408) );
  NAND2_X1 U536 ( .A1(n406), .A2(n390), .ZN(n586) );
  AND2_X2 U537 ( .A1(n408), .A2(n351), .ZN(n407) );
  NAND2_X1 U538 ( .A1(n671), .A2(G234), .ZN(n410) );
  NAND2_X1 U539 ( .A1(n795), .A2(n717), .ZN(n619) );
  NAND2_X1 U540 ( .A1(n416), .A2(n575), .ZN(n577) );
  NAND2_X1 U541 ( .A1(n417), .A2(n514), .ZN(n630) );
  XNOR2_X1 U542 ( .A(n674), .B(n418), .ZN(n787) );
  AND2_X2 U543 ( .A1(n670), .A2(n669), .ZN(n674) );
  INV_X1 U544 ( .A(n593), .ZN(n420) );
  XNOR2_X2 U545 ( .A(n478), .B(G472), .ZN(n593) );
  NAND2_X1 U546 ( .A1(n427), .A2(n371), .ZN(n461) );
  NAND2_X1 U547 ( .A1(n464), .A2(n674), .ZN(n427) );
  XNOR2_X1 U548 ( .A(n449), .B(n656), .ZN(n657) );
  NAND2_X1 U549 ( .A1(n424), .A2(n695), .ZN(n446) );
  XNOR2_X1 U550 ( .A(n426), .B(KEYINPUT72), .ZN(n445) );
  NAND2_X1 U551 ( .A1(n437), .A2(n440), .ZN(n426) );
  OR2_X1 U552 ( .A1(n427), .A2(n369), .ZN(n454) );
  XNOR2_X1 U553 ( .A(n444), .B(n621), .ZN(n672) );
  OR2_X2 U554 ( .A1(n677), .A2(G902), .ZN(n478) );
  XNOR2_X2 U555 ( .A(n512), .B(n511), .ZN(n706) );
  AND2_X2 U556 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U557 ( .A1(n706), .A2(n513), .ZN(n432) );
  AND2_X1 U558 ( .A1(n624), .A2(n434), .ZN(n650) );
  NAND2_X1 U559 ( .A1(n436), .A2(n447), .ZN(n435) );
  XNOR2_X1 U560 ( .A(n590), .B(n448), .ZN(n436) );
  NAND2_X1 U561 ( .A1(n453), .A2(n607), .ZN(n589) );
  XNOR2_X1 U562 ( .A(n439), .B(n438), .ZN(n437) );
  INV_X1 U563 ( .A(KEYINPUT67), .ZN(n438) );
  INV_X1 U564 ( .A(n619), .ZN(n440) );
  NOR2_X2 U565 ( .A1(n676), .A2(n729), .ZN(n699) );
  NAND2_X1 U566 ( .A1(n445), .A2(n620), .ZN(n444) );
  XNOR2_X2 U567 ( .A(n530), .B(n529), .ZN(n648) );
  NAND2_X1 U568 ( .A1(n451), .A2(n450), .ZN(n449) );
  INV_X1 U569 ( .A(n655), .ZN(n450) );
  XNOR2_X2 U570 ( .A(n569), .B(n568), .ZN(n655) );
  XNOR2_X1 U571 ( .A(n452), .B(n654), .ZN(n451) );
  NAND2_X1 U572 ( .A1(n671), .A2(KEYINPUT65), .ZN(n457) );
  INV_X1 U573 ( .A(n671), .ZN(n460) );
  INV_X1 U574 ( .A(n672), .ZN(n464) );
  BUF_X1 U575 ( .A(n699), .Z(n705) );
  XOR2_X1 U576 ( .A(n515), .B(n477), .Z(n465) );
  XOR2_X1 U577 ( .A(KEYINPUT82), .B(n496), .Z(n466) );
  INV_X1 U578 ( .A(KEYINPUT75), .ZN(n654) );
  XNOR2_X1 U579 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U580 ( .A(n522), .B(n521), .ZN(n524) );
  XNOR2_X1 U581 ( .A(n512), .B(n465), .ZN(n677) );
  XNOR2_X2 U582 ( .A(G143), .B(KEYINPUT81), .ZN(n467) );
  XNOR2_X1 U583 ( .A(n468), .B(KEYINPUT69), .ZN(n469) );
  XNOR2_X2 U584 ( .A(n525), .B(n469), .ZN(n786) );
  XNOR2_X2 U585 ( .A(n786), .B(G146), .ZN(n512) );
  XNOR2_X1 U586 ( .A(n471), .B(n470), .ZN(n473) );
  XOR2_X1 U587 ( .A(G101), .B(G113), .Z(n472) );
  NAND2_X1 U588 ( .A1(n550), .A2(G210), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n474), .B(G137), .ZN(n476) );
  XNOR2_X1 U590 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n475) );
  XNOR2_X1 U591 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n481) );
  XOR2_X1 U593 ( .A(KEYINPUT84), .B(G119), .Z(n483) );
  XNOR2_X1 U594 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U595 ( .A(G137), .B(G140), .Z(n505) );
  INV_X1 U596 ( .A(n505), .ZN(n485) );
  NAND2_X1 U597 ( .A1(n700), .A2(n429), .ZN(n489) );
  XOR2_X1 U598 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n486) );
  XNOR2_X2 U599 ( .A(G902), .B(KEYINPUT15), .ZN(n671) );
  XOR2_X1 U600 ( .A(KEYINPUT95), .B(n487), .Z(n488) );
  XNOR2_X1 U601 ( .A(n490), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U602 ( .A1(G952), .A2(n493), .ZN(n491) );
  XNOR2_X1 U603 ( .A(KEYINPUT94), .B(n491), .ZN(n763) );
  NOR2_X1 U604 ( .A1(G953), .A2(n763), .ZN(n572) );
  AND2_X1 U605 ( .A1(G902), .A2(n493), .ZN(n571) );
  NAND2_X1 U606 ( .A1(n492), .A2(n571), .ZN(n494) );
  NOR2_X1 U607 ( .A1(G900), .A2(n494), .ZN(n495) );
  NOR2_X1 U608 ( .A1(n572), .A2(n495), .ZN(n496) );
  NAND2_X1 U609 ( .A1(n497), .A2(G221), .ZN(n499) );
  INV_X1 U610 ( .A(KEYINPUT21), .ZN(n498) );
  XNOR2_X1 U611 ( .A(n499), .B(n498), .ZN(n733) );
  NAND2_X1 U612 ( .A1(n466), .A2(n733), .ZN(n500) );
  XNOR2_X1 U613 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n502) );
  INV_X1 U614 ( .A(KEYINPUT109), .ZN(n501) );
  INV_X1 U615 ( .A(G227), .ZN(n504) );
  OR2_X1 U616 ( .A1(n492), .A2(n504), .ZN(n507) );
  XOR2_X1 U617 ( .A(G101), .B(n505), .Z(n506) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n510) );
  XNOR2_X1 U619 ( .A(n509), .B(n508), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n510), .B(n516), .ZN(n511) );
  INV_X1 U621 ( .A(G469), .ZN(n513) );
  XNOR2_X1 U622 ( .A(G122), .B(n516), .ZN(n517) );
  NAND2_X1 U623 ( .A1(n479), .A2(G224), .ZN(n522) );
  XOR2_X1 U624 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n520) );
  XNOR2_X1 U625 ( .A(n524), .B(n523), .ZN(n527) );
  INV_X1 U626 ( .A(n525), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U628 ( .A1(n685), .A2(n671), .ZN(n530) );
  NAND2_X1 U629 ( .A1(G210), .A2(n531), .ZN(n529) );
  NAND2_X1 U630 ( .A1(G214), .A2(n531), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n532), .B(KEYINPUT93), .ZN(n753) );
  INV_X1 U632 ( .A(n534), .ZN(n719) );
  NAND2_X1 U633 ( .A1(G217), .A2(n535), .ZN(n536) );
  XNOR2_X1 U634 ( .A(n354), .B(n536), .ZN(n543) );
  XNOR2_X1 U635 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U636 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n540) );
  XOR2_X1 U637 ( .A(n541), .B(n540), .Z(n542) );
  INV_X1 U638 ( .A(G478), .ZN(n544) );
  XOR2_X1 U639 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n546) );
  XNOR2_X1 U640 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n545) );
  XNOR2_X1 U641 ( .A(n549), .B(n548), .ZN(n552) );
  AND2_X1 U642 ( .A1(n550), .A2(G214), .ZN(n551) );
  XNOR2_X1 U643 ( .A(n552), .B(n551), .ZN(n556) );
  XNOR2_X1 U644 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U645 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U646 ( .A1(n692), .A2(n429), .ZN(n559) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(G475), .Z(n558) );
  INV_X1 U648 ( .A(n591), .ZN(n599) );
  NOR2_X2 U649 ( .A1(n600), .A2(n599), .ZN(n724) );
  INV_X1 U650 ( .A(n724), .ZN(n560) );
  NOR2_X1 U651 ( .A1(n719), .A2(n560), .ZN(n562) );
  XNOR2_X1 U652 ( .A(G146), .B(KEYINPUT115), .ZN(n561) );
  XNOR2_X1 U653 ( .A(n562), .B(n561), .ZN(G48) );
  INV_X1 U654 ( .A(n753), .ZN(n623) );
  AND2_X1 U655 ( .A1(n724), .A2(n623), .ZN(n563) );
  INV_X1 U656 ( .A(n648), .ZN(n664) );
  XNOR2_X1 U657 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n564) );
  XNOR2_X1 U658 ( .A(n564), .B(KEYINPUT89), .ZN(n565) );
  XNOR2_X1 U659 ( .A(n566), .B(n565), .ZN(n567) );
  INV_X1 U660 ( .A(KEYINPUT112), .ZN(n568) );
  XNOR2_X1 U661 ( .A(G125), .B(KEYINPUT37), .ZN(n570) );
  XNOR2_X1 U662 ( .A(n655), .B(n570), .ZN(G27) );
  INV_X1 U663 ( .A(G953), .ZN(n776) );
  NOR2_X1 U664 ( .A1(G898), .A2(n776), .ZN(n775) );
  NAND2_X1 U665 ( .A1(n775), .A2(n571), .ZN(n574) );
  INV_X1 U666 ( .A(n572), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U668 ( .A(KEYINPUT0), .ZN(n576) );
  XNOR2_X2 U669 ( .A(n577), .B(n576), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n600), .A2(n591), .ZN(n749) );
  AND2_X1 U671 ( .A1(n749), .A2(n733), .ZN(n578) );
  NAND2_X1 U672 ( .A1(n594), .A2(n578), .ZN(n580) );
  INV_X1 U673 ( .A(n586), .ZN(n581) );
  INV_X1 U674 ( .A(n734), .ZN(n611) );
  NOR2_X1 U675 ( .A1(n581), .A2(n611), .ZN(n583) );
  INV_X1 U676 ( .A(n607), .ZN(n582) );
  NAND2_X1 U677 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U678 ( .A1(n610), .A2(n584), .ZN(n602) );
  XOR2_X1 U679 ( .A(G101), .B(n602), .Z(G3) );
  NAND2_X1 U680 ( .A1(n585), .A2(n733), .ZN(n731) );
  XNOR2_X1 U681 ( .A(KEYINPUT91), .B(KEYINPUT33), .ZN(n587) );
  XNOR2_X1 U682 ( .A(n587), .B(KEYINPUT71), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n600), .A2(n591), .ZN(n647) );
  XOR2_X1 U684 ( .A(n592), .B(G122), .Z(G24) );
  NAND2_X1 U685 ( .A1(n592), .A2(KEYINPUT44), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n741), .A2(n596), .ZN(n595) );
  INV_X1 U687 ( .A(n596), .ZN(n598) );
  NOR2_X1 U688 ( .A1(n598), .A2(n597), .ZN(n713) );
  NOR2_X1 U689 ( .A1(n601), .A2(n747), .ZN(n603) );
  NOR2_X1 U690 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U692 ( .A(n606), .B(KEYINPUT88), .ZN(n617) );
  OR2_X1 U693 ( .A1(n586), .A2(n734), .ZN(n608) );
  OR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U695 ( .A(n610), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n586), .A2(n611), .ZN(n613) );
  NOR2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n717) );
  AND2_X1 U699 ( .A1(n619), .A2(KEYINPUT44), .ZN(n616) );
  NOR2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n620) );
  INV_X1 U701 ( .A(KEYINPUT45), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n362), .A2(n466), .ZN(n622) );
  INV_X1 U703 ( .A(KEYINPUT38), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n648), .B(n625), .ZN(n752) );
  INV_X1 U705 ( .A(n752), .ZN(n626) );
  XNOR2_X1 U706 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(KEYINPUT73), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n753), .A2(n752), .ZN(n748) );
  NAND2_X1 U709 ( .A1(n748), .A2(n749), .ZN(n629) );
  XOR2_X1 U710 ( .A(KEYINPUT41), .B(n629), .Z(n764) );
  NOR2_X1 U711 ( .A1(n764), .A2(n630), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT42), .ZN(n797) );
  INV_X1 U713 ( .A(n797), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n635) );
  INV_X1 U715 ( .A(KEYINPUT46), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n635), .B(n634), .ZN(n658) );
  INV_X1 U717 ( .A(KEYINPUT47), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n644), .A2(KEYINPUT76), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n534), .A2(n360), .ZN(n638) );
  INV_X1 U720 ( .A(KEYINPUT83), .ZN(n645) );
  OR2_X1 U721 ( .A1(n747), .A2(n645), .ZN(n637) );
  OR2_X1 U722 ( .A1(n639), .A2(KEYINPUT76), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n747), .A2(n645), .ZN(n643) );
  AND2_X1 U725 ( .A1(KEYINPUT47), .A2(KEYINPUT76), .ZN(n642) );
  AND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  OR2_X1 U727 ( .A1(n364), .A2(n646), .ZN(n651) );
  NOR2_X1 U728 ( .A1(n353), .A2(n647), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n723) );
  NAND2_X1 U730 ( .A1(n651), .A2(n723), .ZN(n652) );
  INV_X1 U731 ( .A(KEYINPUT70), .ZN(n656) );
  INV_X1 U732 ( .A(KEYINPUT48), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n726), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT113), .ZN(n796) );
  NAND2_X1 U735 ( .A1(n365), .A2(n586), .ZN(n663) );
  XOR2_X1 U736 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n665) );
  OR2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n667) );
  INV_X1 U739 ( .A(KEYINPUT107), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n794) );
  INV_X1 U741 ( .A(n794), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n796), .A2(n668), .ZN(n669) );
  BUF_X1 U743 ( .A(n672), .Z(n673) );
  NAND2_X1 U744 ( .A1(n674), .A2(KEYINPUT2), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n673), .A2(n675), .ZN(n729) );
  NAND2_X1 U746 ( .A1(n699), .A2(G472), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n681) );
  INV_X1 U748 ( .A(G952), .ZN(n680) );
  NAND2_X1 U749 ( .A1(n681), .A2(n695), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U751 ( .A1(n699), .A2(G210), .ZN(n687) );
  XNOR2_X1 U752 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n683) );
  XOR2_X1 U753 ( .A(n683), .B(KEYINPUT55), .Z(n684) );
  XNOR2_X1 U754 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n688), .A2(n695), .ZN(n690) );
  XNOR2_X1 U756 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n690), .B(n689), .ZN(G51) );
  INV_X1 U758 ( .A(n695), .ZN(n710) );
  NAND2_X1 U759 ( .A1(n699), .A2(G475), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n691) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n698) );
  INV_X1 U763 ( .A(KEYINPUT60), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n698), .B(n697), .ZN(G60) );
  NAND2_X1 U765 ( .A1(n705), .A2(G217), .ZN(n703) );
  XNOR2_X1 U766 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n700), .B(n701), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U769 ( .A1(n704), .A2(n710), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n705), .A2(G469), .ZN(n709) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  XNOR2_X1 U772 ( .A(n352), .B(n707), .ZN(n708) );
  XNOR2_X1 U773 ( .A(n709), .B(n708), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n713), .A2(n724), .ZN(n712) );
  XNOR2_X1 U776 ( .A(n712), .B(G104), .ZN(G6) );
  XOR2_X1 U777 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n715) );
  NAND2_X1 U778 ( .A1(n713), .A2(n726), .ZN(n714) );
  XNOR2_X1 U779 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U780 ( .A(G107), .B(n716), .ZN(G9) );
  XNOR2_X1 U781 ( .A(G110), .B(n717), .ZN(G12) );
  INV_X1 U782 ( .A(n726), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U784 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n720) );
  XNOR2_X1 U785 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U786 ( .A(G128), .B(n722), .ZN(G30) );
  XNOR2_X1 U787 ( .A(G143), .B(n723), .ZN(G45) );
  NAND2_X1 U788 ( .A1(n724), .A2(n727), .ZN(n725) );
  XNOR2_X1 U789 ( .A(G113), .B(n725), .ZN(G15) );
  NAND2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U791 ( .A(n728), .B(G116), .ZN(G18) );
  NOR2_X1 U792 ( .A1(n359), .A2(n729), .ZN(n730) );
  XNOR2_X1 U793 ( .A(n730), .B(KEYINPUT85), .ZN(n771) );
  NAND2_X1 U794 ( .A1(n586), .A2(n731), .ZN(n732) );
  XOR2_X1 U795 ( .A(KEYINPUT50), .B(n732), .Z(n738) );
  NOR2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U797 ( .A(n735), .B(KEYINPUT49), .ZN(n736) );
  NOR2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U799 ( .A(n739), .B(KEYINPUT116), .ZN(n740) );
  NOR2_X1 U800 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U801 ( .A(KEYINPUT51), .B(n742), .Z(n743) );
  NOR2_X1 U802 ( .A1(n764), .A2(n743), .ZN(n744) );
  XOR2_X1 U803 ( .A(KEYINPUT117), .B(n744), .Z(n760) );
  BUF_X1 U804 ( .A(n745), .Z(n746) );
  INV_X1 U805 ( .A(n746), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n748), .A2(n379), .ZN(n751) );
  INV_X1 U807 ( .A(n749), .ZN(n750) );
  NAND2_X1 U808 ( .A1(n751), .A2(n750), .ZN(n755) );
  NAND2_X1 U809 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U810 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U812 ( .A(n758), .B(KEYINPUT118), .ZN(n759) );
  NOR2_X1 U813 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U814 ( .A(n761), .B(KEYINPUT52), .ZN(n762) );
  NOR2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n768) );
  INV_X1 U816 ( .A(n764), .ZN(n765) );
  NAND2_X1 U817 ( .A1(n746), .A2(n765), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n766), .B(KEYINPUT119), .ZN(n767) );
  NOR2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U820 ( .A(KEYINPUT120), .B(n769), .ZN(n770) );
  NAND2_X1 U821 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U822 ( .A1(n772), .A2(G953), .ZN(n773) );
  XNOR2_X1 U823 ( .A(n773), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U824 ( .A1(n775), .A2(n774), .ZN(n784) );
  INV_X1 U825 ( .A(n673), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U827 ( .A1(G953), .A2(G224), .ZN(n778) );
  XNOR2_X1 U828 ( .A(KEYINPUT61), .B(n778), .ZN(n779) );
  NAND2_X1 U829 ( .A1(n779), .A2(G898), .ZN(n780) );
  NAND2_X1 U830 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U831 ( .A(n782), .B(KEYINPUT126), .ZN(n783) );
  XNOR2_X1 U832 ( .A(n784), .B(n783), .ZN(G69) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(n788) );
  NAND2_X1 U834 ( .A1(n787), .A2(n479), .ZN(n793) );
  XNOR2_X1 U835 ( .A(n788), .B(G227), .ZN(n789) );
  NAND2_X1 U836 ( .A1(n789), .A2(G900), .ZN(n790) );
  XOR2_X1 U837 ( .A(KEYINPUT127), .B(n790), .Z(n791) );
  NAND2_X1 U838 ( .A1(n791), .A2(G953), .ZN(n792) );
  NAND2_X1 U839 ( .A1(n793), .A2(n792), .ZN(G72) );
  XNOR2_X1 U840 ( .A(G140), .B(n794), .ZN(G42) );
  XNOR2_X1 U841 ( .A(G119), .B(n795), .ZN(G21) );
  XOR2_X1 U842 ( .A(G134), .B(n796), .Z(G36) );
  XOR2_X1 U843 ( .A(G137), .B(n797), .Z(G39) );
endmodule

