

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n526), .B(n525), .ZN(n900) );
  AND2_X1 U556 ( .A1(n527), .A2(G2104), .ZN(n899) );
  NOR2_X1 U557 ( .A1(n667), .A2(n957), .ZN(n615) );
  OR2_X1 U558 ( .A1(n624), .A2(n990), .ZN(n626) );
  OR2_X1 U559 ( .A1(n666), .A2(n665), .ZN(n682) );
  NOR2_X1 U560 ( .A1(G651), .A2(n578), .ZN(n791) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n798) );
  NAND2_X1 U562 ( .A1(n900), .A2(G138), .ZN(n529) );
  XNOR2_X1 U563 ( .A(n533), .B(KEYINPUT23), .ZN(n534) );
  INV_X1 U564 ( .A(KEYINPUT64), .ZN(n533) );
  OR2_X1 U565 ( .A1(n711), .A2(n710), .ZN(n521) );
  AND2_X1 U566 ( .A1(n987), .A2(n756), .ZN(n522) );
  INV_X1 U567 ( .A(KEYINPUT26), .ZN(n614) );
  NOR2_X1 U568 ( .A1(n993), .A2(n618), .ZN(n624) );
  INV_X1 U569 ( .A(KEYINPUT97), .ZN(n625) );
  XNOR2_X1 U570 ( .A(KEYINPUT98), .B(KEYINPUT30), .ZN(n656) );
  XNOR2_X1 U571 ( .A(n657), .B(n656), .ZN(n658) );
  AND2_X1 U572 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U573 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U574 ( .A1(n652), .A2(n651), .ZN(n675) );
  INV_X1 U575 ( .A(KEYINPUT100), .ZN(n692) );
  XNOR2_X1 U576 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U577 ( .A(KEYINPUT70), .B(KEYINPUT13), .ZN(n608) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n743), .A2(n522), .ZN(n744) );
  XNOR2_X1 U580 ( .A(n609), .B(n608), .ZN(n610) );
  NOR2_X1 U581 ( .A1(n578), .A2(n545), .ZN(n795) );
  XNOR2_X1 U582 ( .A(n535), .B(n534), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n613), .A2(n612), .ZN(n993) );
  NOR2_X1 U584 ( .A1(n541), .A2(n540), .ZN(G160) );
  INV_X1 U585 ( .A(G2105), .ZN(n527) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n902) );
  NAND2_X1 U587 ( .A1(G114), .A2(n902), .ZN(n524) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n527), .ZN(n903) );
  NAND2_X1 U589 ( .A1(G126), .A2(n903), .ZN(n523) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n532) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  NAND2_X1 U592 ( .A1(G102), .A2(n899), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT89), .B(n530), .Z(n531) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G101), .A2(n899), .ZN(n535) );
  NAND2_X1 U597 ( .A1(G137), .A2(n900), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G113), .A2(n902), .ZN(n539) );
  NAND2_X1 U600 ( .A1(G125), .A2(n903), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U602 ( .A(G543), .B(KEYINPUT0), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n542), .B(KEYINPUT65), .ZN(n578) );
  INV_X1 U604 ( .A(G651), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G75), .A2(n795), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G88), .A2(n798), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n550) );
  NOR2_X1 U608 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT1), .B(n546), .Z(n789) );
  NAND2_X1 U610 ( .A1(G62), .A2(n789), .ZN(n548) );
  NAND2_X1 U611 ( .A1(G50), .A2(n791), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U613 ( .A1(n550), .A2(n549), .ZN(G166) );
  INV_X1 U614 ( .A(G166), .ZN(G303) );
  NAND2_X1 U615 ( .A1(n791), .A2(G52), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n789), .A2(G64), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G77), .A2(n795), .ZN(n554) );
  NAND2_X1 U619 ( .A1(G90), .A2(n798), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G63), .A2(n789), .ZN(n559) );
  NAND2_X1 U625 ( .A1(G51), .A2(n791), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT6), .B(n560), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n798), .A2(G89), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G76), .A2(n795), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U632 ( .A(n564), .B(KEYINPUT5), .Z(n565) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT74), .B(n567), .Z(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT7), .B(n568), .ZN(G168) );
  XNOR2_X1 U636 ( .A(KEYINPUT75), .B(KEYINPUT8), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(G168), .ZN(G286) );
  NAND2_X1 U638 ( .A1(G48), .A2(n791), .ZN(n576) );
  NAND2_X1 U639 ( .A1(G86), .A2(n798), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G61), .A2(n789), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n795), .A2(G73), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n572), .Z(n573) );
  NOR2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U647 ( .A1(G49), .A2(n791), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G87), .A2(n578), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U650 ( .A1(n789), .A2(n581), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G651), .A2(G74), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(G288) );
  NAND2_X1 U653 ( .A1(G72), .A2(n795), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G60), .A2(n789), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G85), .A2(n798), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G47), .A2(n791), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  OR2_X1 U659 ( .A1(n589), .A2(n588), .ZN(G290) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n730) );
  INV_X1 U661 ( .A(n730), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G160), .A2(G40), .ZN(n729) );
  OR2_X2 U663 ( .A1(n590), .A2(n729), .ZN(n667) );
  NAND2_X1 U664 ( .A1(n667), .A2(G8), .ZN(n695) );
  NOR2_X1 U665 ( .A1(G2090), .A2(G303), .ZN(n591) );
  XNOR2_X1 U666 ( .A(KEYINPUT102), .B(n591), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n592), .A2(G8), .ZN(n683) );
  NAND2_X1 U668 ( .A1(G92), .A2(n798), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G66), .A2(n789), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U671 ( .A(n595), .B(KEYINPUT71), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G79), .A2(n795), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G54), .A2(n791), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U675 ( .A(KEYINPUT72), .B(n598), .Z(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT15), .ZN(n990) );
  XOR2_X1 U678 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n603) );
  NAND2_X1 U679 ( .A1(G56), .A2(n789), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n603), .B(n602), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n795), .A2(G68), .ZN(n604) );
  XNOR2_X1 U682 ( .A(KEYINPUT69), .B(n604), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n798), .A2(G81), .ZN(n605) );
  XOR2_X1 U684 ( .A(n605), .B(KEYINPUT12), .Z(n606) );
  NOR2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n791), .A2(G43), .ZN(n612) );
  INV_X1 U688 ( .A(G1996), .ZN(n957) );
  XNOR2_X1 U689 ( .A(n615), .B(n614), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n667), .A2(G1341), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n990), .A2(n624), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT96), .B(n619), .ZN(n623) );
  NOR2_X1 U694 ( .A1(G2067), .A2(n667), .ZN(n621) );
  INV_X1 U695 ( .A(n667), .ZN(n648) );
  NOR2_X1 U696 ( .A1(n648), .A2(G1348), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n640) );
  XNOR2_X1 U699 ( .A(n626), .B(n625), .ZN(n638) );
  NAND2_X1 U700 ( .A1(G65), .A2(n789), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G53), .A2(n791), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G78), .A2(n795), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G91), .A2(n798), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n805) );
  NAND2_X1 U707 ( .A1(n648), .A2(G2072), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT27), .ZN(n635) );
  AND2_X1 U709 ( .A1(G1956), .A2(n667), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n642) );
  NOR2_X1 U711 ( .A1(n805), .A2(n642), .ZN(n637) );
  INV_X1 U712 ( .A(KEYINPUT28), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n641) );
  AND2_X1 U714 ( .A1(n638), .A2(n641), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n646) );
  INV_X1 U716 ( .A(n641), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n805), .A2(n642), .ZN(n643) );
  OR2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U719 ( .A(KEYINPUT29), .B(n647), .Z(n652) );
  NAND2_X1 U720 ( .A1(G1961), .A2(n667), .ZN(n650) );
  XOR2_X1 U721 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NAND2_X1 U722 ( .A1(n648), .A2(n961), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n653) );
  OR2_X1 U724 ( .A1(G301), .A2(n653), .ZN(n651) );
  NAND2_X1 U725 ( .A1(G301), .A2(n653), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(KEYINPUT99), .ZN(n660) );
  NOR2_X1 U727 ( .A1(G1966), .A2(n695), .ZN(n663) );
  NOR2_X1 U728 ( .A1(G2084), .A2(n667), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G8), .A2(n655), .ZN(n657) );
  NOR2_X1 U731 ( .A1(G168), .A2(n658), .ZN(n659) );
  XOR2_X1 U732 ( .A(KEYINPUT31), .B(n661), .Z(n673) );
  AND2_X1 U733 ( .A1(n675), .A2(n673), .ZN(n666) );
  AND2_X1 U734 ( .A1(G8), .A2(n662), .ZN(n664) );
  OR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  INV_X1 U736 ( .A(G8), .ZN(n672) );
  NOR2_X1 U737 ( .A1(G1971), .A2(n695), .ZN(n669) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(G303), .ZN(n671) );
  OR2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U742 ( .A1(n673), .A2(n676), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n679) );
  INV_X1 U744 ( .A(n676), .ZN(n677) );
  OR2_X1 U745 ( .A1(n677), .A2(G286), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT32), .ZN(n681) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n691) );
  NAND2_X1 U749 ( .A1(n683), .A2(n691), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n695), .A2(n684), .ZN(n689) );
  INV_X1 U751 ( .A(n695), .ZN(n697) );
  NOR2_X1 U752 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XOR2_X1 U753 ( .A(n685), .B(KEYINPUT24), .Z(n686) );
  XNOR2_X1 U754 ( .A(KEYINPUT95), .B(n686), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n697), .A2(n687), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n711) );
  NOR2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n696) );
  NOR2_X1 U758 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n696), .A2(n690), .ZN(n982) );
  NAND2_X1 U760 ( .A1(n691), .A2(n982), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n703) );
  NAND2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U763 ( .A(KEYINPUT33), .ZN(n705) );
  NAND2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U765 ( .A1(n705), .A2(n698), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT101), .ZN(n704) );
  AND2_X1 U767 ( .A1(n981), .A2(n704), .ZN(n701) );
  XNOR2_X1 U768 ( .A(G1981), .B(G305), .ZN(n995) );
  INV_X1 U769 ( .A(n995), .ZN(n700) );
  AND2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n709) );
  INV_X1 U772 ( .A(n704), .ZN(n706) );
  OR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  OR2_X1 U774 ( .A1(n995), .A2(n707), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U776 ( .A1(G95), .A2(n899), .ZN(n712) );
  XNOR2_X1 U777 ( .A(n712), .B(KEYINPUT92), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G119), .A2(n903), .ZN(n713) );
  XOR2_X1 U779 ( .A(KEYINPUT91), .B(n713), .Z(n714) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U781 ( .A1(G107), .A2(n902), .ZN(n717) );
  NAND2_X1 U782 ( .A1(G131), .A2(n900), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n896) );
  XOR2_X1 U785 ( .A(KEYINPUT93), .B(G1991), .Z(n962) );
  AND2_X1 U786 ( .A1(n896), .A2(n962), .ZN(n728) );
  NAND2_X1 U787 ( .A1(G117), .A2(n902), .ZN(n721) );
  NAND2_X1 U788 ( .A1(G129), .A2(n903), .ZN(n720) );
  NAND2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U790 ( .A1(n899), .A2(G105), .ZN(n722) );
  XOR2_X1 U791 ( .A(KEYINPUT38), .B(n722), .Z(n723) );
  NOR2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U793 ( .A1(n900), .A2(G141), .ZN(n725) );
  NAND2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n895) );
  AND2_X1 U795 ( .A1(n895), .A2(G1996), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n939) );
  NOR2_X1 U797 ( .A1(n730), .A2(n729), .ZN(n756) );
  XOR2_X1 U798 ( .A(KEYINPUT94), .B(n756), .Z(n731) );
  NOR2_X1 U799 ( .A1(n939), .A2(n731), .ZN(n748) );
  INV_X1 U800 ( .A(n748), .ZN(n742) );
  XNOR2_X1 U801 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n735) );
  NAND2_X1 U802 ( .A1(G104), .A2(n899), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G140), .A2(n900), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U805 ( .A(n735), .B(n734), .ZN(n740) );
  NAND2_X1 U806 ( .A1(G116), .A2(n902), .ZN(n737) );
  NAND2_X1 U807 ( .A1(G128), .A2(n903), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U809 ( .A(KEYINPUT35), .B(n738), .Z(n739) );
  NOR2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U811 ( .A(KEYINPUT36), .B(n741), .ZN(n917) );
  XNOR2_X1 U812 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NOR2_X1 U813 ( .A1(n917), .A2(n753), .ZN(n949) );
  NAND2_X1 U814 ( .A1(n756), .A2(n949), .ZN(n751) );
  NAND2_X1 U815 ( .A1(n742), .A2(n751), .ZN(n743) );
  XNOR2_X1 U816 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U817 ( .A1(n521), .A2(n744), .ZN(n759) );
  NOR2_X1 U818 ( .A1(G1996), .A2(n895), .ZN(n929) );
  NOR2_X1 U819 ( .A1(n962), .A2(n896), .ZN(n932) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n745) );
  XOR2_X1 U821 ( .A(n745), .B(KEYINPUT103), .Z(n746) );
  NOR2_X1 U822 ( .A1(n932), .A2(n746), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U824 ( .A1(n929), .A2(n749), .ZN(n750) );
  XNOR2_X1 U825 ( .A(KEYINPUT39), .B(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n917), .A2(n753), .ZN(n933) );
  NAND2_X1 U828 ( .A1(n754), .A2(n933), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U830 ( .A(KEYINPUT104), .B(n757), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U832 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G108), .ZN(G238) );
  INV_X1 U835 ( .A(n805), .ZN(G299) );
  NAND2_X1 U836 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U837 ( .A(n761), .B(KEYINPUT10), .ZN(n762) );
  XNOR2_X1 U838 ( .A(KEYINPUT66), .B(n762), .ZN(G223) );
  INV_X1 U839 ( .A(G223), .ZN(n833) );
  NAND2_X1 U840 ( .A1(n833), .A2(G567), .ZN(n763) );
  XNOR2_X1 U841 ( .A(n763), .B(KEYINPUT67), .ZN(n764) );
  XNOR2_X1 U842 ( .A(KEYINPUT11), .B(n764), .ZN(G234) );
  INV_X1 U843 ( .A(G860), .ZN(n788) );
  OR2_X1 U844 ( .A1(n993), .A2(n788), .ZN(G153) );
  NAND2_X1 U845 ( .A1(G868), .A2(G171), .ZN(n766) );
  INV_X1 U846 ( .A(G868), .ZN(n813) );
  NAND2_X1 U847 ( .A1(n990), .A2(n813), .ZN(n765) );
  NAND2_X1 U848 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U849 ( .A(n767), .B(KEYINPUT73), .ZN(G284) );
  NOR2_X1 U850 ( .A1(G286), .A2(n813), .ZN(n769) );
  NOR2_X1 U851 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U852 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U853 ( .A(KEYINPUT76), .B(n770), .ZN(G297) );
  NAND2_X1 U854 ( .A1(G559), .A2(n788), .ZN(n771) );
  XOR2_X1 U855 ( .A(KEYINPUT77), .B(n771), .Z(n772) );
  NAND2_X1 U856 ( .A1(n772), .A2(n990), .ZN(n773) );
  XNOR2_X1 U857 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(G868), .A2(n993), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G868), .A2(n990), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G559), .A2(n774), .ZN(n775) );
  NOR2_X1 U861 ( .A1(n776), .A2(n775), .ZN(G282) );
  NAND2_X1 U862 ( .A1(G99), .A2(n899), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G111), .A2(n902), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U865 ( .A(KEYINPUT78), .B(n779), .ZN(n784) );
  NAND2_X1 U866 ( .A1(G123), .A2(n903), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT18), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n900), .A2(G135), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n931) );
  XNOR2_X1 U871 ( .A(n931), .B(G2096), .ZN(n786) );
  INV_X1 U872 ( .A(G2100), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(G156) );
  NAND2_X1 U874 ( .A1(G559), .A2(n990), .ZN(n787) );
  XOR2_X1 U875 ( .A(n993), .B(n787), .Z(n810) );
  NAND2_X1 U876 ( .A1(n788), .A2(n810), .ZN(n802) );
  NAND2_X1 U877 ( .A1(n789), .A2(G67), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n790), .B(KEYINPUT80), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U881 ( .A(n794), .B(KEYINPUT81), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G80), .A2(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G93), .A2(n798), .ZN(n799) );
  XNOR2_X1 U885 ( .A(KEYINPUT79), .B(n799), .ZN(n800) );
  NOR2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n812) );
  XOR2_X1 U887 ( .A(n802), .B(n812), .Z(G145) );
  XNOR2_X1 U888 ( .A(G305), .B(n812), .ZN(n809) );
  XOR2_X1 U889 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n803) );
  XNOR2_X1 U890 ( .A(G288), .B(n803), .ZN(n804) );
  XNOR2_X1 U891 ( .A(G290), .B(n804), .ZN(n807) );
  XNOR2_X1 U892 ( .A(n805), .B(G166), .ZN(n806) );
  XNOR2_X1 U893 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n809), .B(n808), .ZN(n849) );
  XOR2_X1 U895 ( .A(n849), .B(n810), .Z(n811) );
  NOR2_X1 U896 ( .A1(n813), .A2(n811), .ZN(n815) );
  AND2_X1 U897 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U898 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U903 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n820) );
  XOR2_X1 U906 ( .A(KEYINPUT87), .B(n820), .Z(n821) );
  NOR2_X1 U907 ( .A1(G238), .A2(n821), .ZN(n822) );
  NAND2_X1 U908 ( .A1(G57), .A2(n822), .ZN(n838) );
  NAND2_X1 U909 ( .A1(n838), .A2(G567), .ZN(n830) );
  XOR2_X1 U910 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n824) );
  NAND2_X1 U911 ( .A1(G132), .A2(G82), .ZN(n823) );
  XNOR2_X1 U912 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U913 ( .A1(n825), .A2(G96), .ZN(n826) );
  NOR2_X1 U914 ( .A1(n826), .A2(G218), .ZN(n827) );
  XNOR2_X1 U915 ( .A(n827), .B(KEYINPUT85), .ZN(n837) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n837), .ZN(n828) );
  XNOR2_X1 U917 ( .A(KEYINPUT86), .B(n828), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n927) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n831) );
  XNOR2_X1 U920 ( .A(KEYINPUT88), .B(n831), .ZN(n832) );
  NOR2_X1 U921 ( .A1(n927), .A2(n832), .ZN(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U925 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  INV_X1 U930 ( .A(G132), .ZN(G219) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G82), .ZN(G220) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U936 ( .A(G1341), .B(G2454), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(G2430), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(G1348), .ZN(n846) );
  XOR2_X1 U939 ( .A(G2443), .B(G2427), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2438), .B(G2446), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U942 ( .A(G2451), .B(G2435), .Z(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n847), .A2(G14), .ZN(n848) );
  XOR2_X1 U946 ( .A(KEYINPUT105), .B(n848), .Z(n922) );
  XOR2_X1 U947 ( .A(KEYINPUT106), .B(n922), .Z(G401) );
  XOR2_X1 U948 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n851) );
  XNOR2_X1 U949 ( .A(G171), .B(n849), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n990), .B(n852), .Z(n853) );
  XNOR2_X1 U952 ( .A(n993), .B(n853), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n854), .B(G286), .ZN(n855) );
  NOR2_X1 U954 ( .A1(G37), .A2(n855), .ZN(G397) );
  XOR2_X1 U955 ( .A(G2100), .B(G2096), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(G2678), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2090), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G227) );
  XNOR2_X1 U964 ( .A(G1976), .B(G2474), .ZN(n873) );
  XOR2_X1 U965 ( .A(G1986), .B(G1971), .Z(n865) );
  XNOR2_X1 U966 ( .A(G1961), .B(G1956), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U968 ( .A(G1991), .B(G1981), .Z(n867) );
  XNOR2_X1 U969 ( .A(G1966), .B(G1996), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U975 ( .A1(G124), .A2(n903), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n874), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G112), .A2(n902), .ZN(n875) );
  XOR2_X1 U978 ( .A(KEYINPUT109), .B(n875), .Z(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G100), .A2(n899), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G136), .A2(n900), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U984 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G106), .A2(n899), .ZN(n883) );
  NAND2_X1 U986 ( .A1(G142), .A2(n900), .ZN(n882) );
  NAND2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n884), .B(KEYINPUT45), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n902), .A2(G118), .ZN(n887) );
  XNOR2_X1 U991 ( .A(n887), .B(KEYINPUT110), .ZN(n889) );
  NAND2_X1 U992 ( .A1(G130), .A2(n903), .ZN(n888) );
  NAND2_X1 U993 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n893) );
  XNOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n892) );
  XNOR2_X1 U996 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U997 ( .A(G162), .B(n894), .ZN(n916) );
  XOR2_X1 U998 ( .A(G164), .B(n895), .Z(n897) );
  XOR2_X1 U999 ( .A(n897), .B(n896), .Z(n898) );
  XOR2_X1 U1000 ( .A(n898), .B(n931), .Z(n914) );
  NAND2_X1 U1001 ( .A1(G103), .A2(n899), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(n900), .A2(G139), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(KEYINPUT113), .B(n901), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(G115), .A2(n902), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(G127), .A2(n903), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1007 ( .A(KEYINPUT47), .B(n906), .Z(n907) );
  XNOR2_X1 U1008 ( .A(KEYINPUT114), .B(n907), .ZN(n908) );
  NOR2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n912), .B(KEYINPUT115), .ZN(n940) );
  XNOR2_X1 U1012 ( .A(G160), .B(n940), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1015 ( .A(n918), .B(n917), .Z(n919) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n919), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n920) );
  XOR2_X1 U1018 ( .A(KEYINPUT118), .B(n920), .Z(n921) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G397), .A2(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G395), .A2(n927), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n927), .ZN(G319) );
  INV_X1 U1026 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n930), .Z(n947) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G160), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(KEYINPUT119), .B(n935), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1036 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n950), .ZN(n951) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n974) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n974), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(G29), .ZN(n1034) );
  XOR2_X1 U1047 ( .A(KEYINPUT121), .B(G34), .Z(n954) );
  XNOR2_X1 U1048 ( .A(G2084), .B(KEYINPUT54), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n954), .B(n953), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G35), .B(G2090), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n972) );
  XNOR2_X1 U1052 ( .A(G32), .B(n957), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n961), .B(G27), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G25), .B(n962), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1062 ( .A(n969), .B(KEYINPUT53), .Z(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT120), .B(n970), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1066 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n977), .ZN(n1032) );
  INV_X1 U1069 ( .A(G16), .ZN(n1028) );
  XOR2_X1 U1070 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n978) );
  XNOR2_X1 U1071 ( .A(n1028), .B(n978), .ZN(n1003) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G299), .B(G1956), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n984) );
  AND2_X1 U1076 ( .A1(G303), .A2(G1971), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT124), .B(n985), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1081 ( .A(G1348), .B(n990), .Z(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n1001) );
  XNOR2_X1 U1083 ( .A(n993), .B(G1341), .ZN(n999) );
  XOR2_X1 U1084 ( .A(G168), .B(G1966), .Z(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1086 ( .A(KEYINPUT123), .B(n996), .Z(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT57), .B(n997), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1030) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(n1004), .B(G4), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G6), .B(G1981), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(KEYINPUT125), .B(G1956), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(G20), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1012), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G5), .B(G1961), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1025) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1021) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G1976), .B(G23), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(n1019), .B(KEYINPUT126), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1022), .Z(n1023) );
  XNOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

