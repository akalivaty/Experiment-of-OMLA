//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT93), .B1(new_n202), .B2(G57gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT93), .ZN(new_n204));
  INV_X1    g003(.A(G57gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(G64gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n206), .C1(new_n205), .C2(G64gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT9), .ZN(new_n209));
  NOR2_X1   g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n209), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(new_n210), .ZN(new_n212));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT94), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n211), .A2(KEYINPUT94), .A3(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT21), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G1gat), .B2(new_n222), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(G8gat), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n221), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(G231gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n228), .B2(new_n230), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G155gat), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n236), .B(KEYINPUT95), .Z(new_n237));
  NOR3_X1   g036(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n228), .A2(new_n230), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n231), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n241), .B2(new_n233), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n220), .A2(KEYINPUT21), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G211gat), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n243), .B(new_n245), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n238), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n237), .B1(new_n234), .B2(new_n235), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n241), .A2(new_n233), .A3(new_n239), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT7), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT7), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G85gat), .A3(G92gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n254), .A2(new_n256), .B1(KEYINPUT8), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT96), .B(G92gat), .ZN(new_n259));
  INV_X1    g058(.A(G85gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G99gat), .B(G106gat), .Z(new_n262));
  AND3_X1   g061(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n258), .B2(new_n261), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT89), .ZN(new_n266));
  INV_X1    g065(.A(G43gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G50gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT15), .B1(new_n268), .B2(KEYINPUT87), .ZN(new_n269));
  INV_X1    g068(.A(G50gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G43gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n271), .B(new_n268), .C1(KEYINPUT87), .C2(KEYINPUT15), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT14), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G29gat), .B2(G36gat), .ZN(new_n277));
  INV_X1    g076(.A(G29gat), .ZN(new_n278));
  INV_X1    g077(.A(G36gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT14), .ZN(new_n280));
  NAND2_X1  g079(.A1(G29gat), .A2(G36gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT88), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT88), .B1(G29gat), .B2(G36gat), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n277), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n266), .B1(new_n275), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(KEYINPUT89), .A3(new_n274), .A4(new_n273), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n272), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(new_n277), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n281), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT15), .B(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT17), .B1(new_n296), .B2(KEYINPUT90), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299));
  AOI211_X1 g098(.A(new_n298), .B(new_n299), .C1(new_n289), .C2(new_n295), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n265), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n265), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G190gat), .B(G218gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n301), .A2(new_n308), .A3(new_n302), .A4(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n313), .A3(new_n309), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n252), .A2(new_n317), .A3(KEYINPUT97), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT97), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n247), .B1(new_n238), .B2(new_n242), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n249), .A2(new_n250), .A3(new_n246), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n315), .A2(new_n316), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n326));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G183gat), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT28), .B1(new_n331), .B2(KEYINPUT65), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT27), .B(G183gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n332), .B(new_n333), .C1(KEYINPUT65), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n229), .A2(KEYINPUT27), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n338), .A3(new_n333), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n339), .B2(KEYINPUT28), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341));
  INV_X1    g140(.A(G169gat), .ZN(new_n342));
  INV_X1    g141(.A(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n335), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT64), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT64), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n361), .A2(G169gat), .A3(G176gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n345), .A2(KEYINPUT23), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(new_n360), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n365), .ZN(new_n368));
  INV_X1    g167(.A(new_n362), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n350), .A2(new_n357), .A3(new_n351), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT25), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT73), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(KEYINPUT29), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  INV_X1    g177(.A(G211gat), .ZN(new_n379));
  INV_X1    g178(.A(G218gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT71), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n384), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(new_n387), .A3(new_n383), .A4(new_n385), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n388), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n354), .B(new_n349), .C1(G183gat), .C2(G190gat), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n360), .B1(new_n366), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n331), .A2(new_n338), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT65), .ZN(new_n400));
  AOI21_X1  g199(.A(G190gat), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n401), .B2(new_n332), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n402), .B2(new_n340), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n367), .A3(new_n375), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n377), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n395), .B1(new_n377), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n329), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n377), .A2(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n394), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n377), .A2(new_n395), .A3(new_n404), .ZN(new_n410));
  INV_X1    g209(.A(new_n329), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n412), .A3(KEYINPUT30), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n405), .A2(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n411), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G148gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G141gat), .ZN(new_n419));
  INV_X1    g218(.A(G141gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G148gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G155gat), .B(G162gat), .ZN(new_n423));
  AND2_X1   g222(.A1(KEYINPUT74), .A2(G162gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT74), .A2(G162gat), .ZN(new_n425));
  INV_X1    g224(.A(G155gat), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT2), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n422), .B(new_n423), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n423), .ZN(new_n430));
  XNOR2_X1  g229(.A(G141gat), .B(G148gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(KEYINPUT2), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n435));
  OAI21_X1  g234(.A(G113gat), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G113gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G120gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440));
  INV_X1    g239(.A(G134gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G127gat), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n441), .A2(G127gat), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n437), .A2(G120gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n437), .A2(G120gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n450));
  OAI211_X1 g249(.A(KEYINPUT67), .B(G134gat), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n441), .B1(new_n452), .B2(new_n448), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n442), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n447), .B(new_n451), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n433), .A2(KEYINPUT3), .B1(new_n444), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n423), .B1(new_n428), .B2(new_n422), .ZN(new_n459));
  OR2_X1    g258(.A1(KEYINPUT74), .A2(G162gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(KEYINPUT74), .A2(G162gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(G155gat), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n431), .B1(new_n462), .B2(KEYINPUT2), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n463), .B2(new_n423), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g265(.A1(new_n458), .A2(new_n429), .A3(new_n465), .A4(new_n432), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n457), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n444), .A2(new_n456), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT4), .B1(new_n469), .B2(new_n433), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n464), .A2(new_n471), .A3(new_n456), .A4(new_n444), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(KEYINPUT5), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n468), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n468), .A2(new_n473), .A3(KEYINPUT79), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT76), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n470), .A2(new_n482), .A3(new_n472), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n456), .A3(new_n444), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n483), .A2(new_n468), .A3(new_n474), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n433), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n474), .B1(new_n487), .B2(new_n484), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT77), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n469), .A2(new_n433), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n444), .A2(new_n456), .B1(new_n429), .B2(new_n432), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n475), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT77), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT5), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n486), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G57gat), .B(G85gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G1gat), .B(G29gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g303(.A(new_n502), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n505), .A3(new_n496), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n497), .A2(KEYINPUT6), .A3(new_n502), .ZN(new_n508));
  AOI211_X1 g307(.A(new_n326), .B(new_n417), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT69), .B1(new_n373), .B2(new_n469), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n444), .A2(new_n456), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT69), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n403), .A2(new_n511), .A3(new_n512), .A4(new_n367), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n373), .A2(new_n469), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n510), .A2(new_n513), .A3(new_n517), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT34), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n520), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT32), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G71gat), .B(G99gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n526), .B1(new_n519), .B2(new_n520), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT70), .B1(new_n535), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT32), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n525), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n538), .B(new_n539), .C1(new_n519), .C2(new_n520), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n523), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  AOI211_X1 g341(.A(new_n540), .B(new_n522), .C1(new_n534), .C2(new_n536), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G50gat), .Z(new_n544));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(G22gat), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n465), .B1(new_n394), .B2(KEYINPUT29), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n433), .ZN(new_n551));
  INV_X1    g350(.A(G228gat), .ZN(new_n552));
  INV_X1    g351(.A(G233gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT75), .B1(new_n433), .B2(KEYINPUT3), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n464), .A2(new_n458), .A3(new_n465), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT29), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n555), .B1(new_n559), .B2(new_n394), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n466), .B2(new_n467), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n389), .A2(new_n391), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n465), .B1(new_n563), .B2(KEYINPUT29), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n562), .A2(new_n394), .B1(new_n564), .B2(new_n433), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n565), .A2(new_n554), .B1(KEYINPUT81), .B2(new_n546), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n549), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n558), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n570), .A3(new_n394), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n554), .A3(new_n551), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n564), .A2(new_n433), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n395), .B2(new_n558), .ZN(new_n575));
  INV_X1    g374(.A(new_n554), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n577), .A3(new_n548), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n542), .A2(new_n543), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n509), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n413), .A2(new_n416), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n506), .A2(new_n504), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n505), .B1(new_n481), .B2(new_n496), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n508), .ZN(new_n587));
  OAI211_X1 g386(.A(KEYINPUT85), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n529), .B1(new_n528), .B2(new_n533), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n535), .A2(KEYINPUT70), .A3(new_n532), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n541), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n522), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n537), .A2(new_n523), .A3(new_n541), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n572), .A2(new_n577), .A3(new_n548), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n548), .B1(new_n572), .B2(new_n577), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT35), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT83), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n487), .A2(new_n484), .A3(new_n474), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n468), .A2(new_n473), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT39), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n468), .B2(new_n473), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n502), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n601), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n583), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT83), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n585), .B1(new_n612), .B2(KEYINPUT40), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n579), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n411), .B1(new_n414), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n615), .B2(new_n414), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n412), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n414), .A2(KEYINPUT84), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT37), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n618), .B(new_n616), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n507), .A2(new_n620), .A3(new_n624), .A4(new_n508), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n614), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n542), .B2(new_n543), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n592), .A2(KEYINPUT36), .A3(new_n593), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n579), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n626), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n599), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n218), .A2(new_n265), .A3(new_n219), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n258), .A2(new_n261), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n262), .A2(KEYINPUT98), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n215), .A3(new_n211), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n303), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n635), .B1(new_n637), .B2(new_n641), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n647), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n226), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n291), .B(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n272), .B1(new_n654), .B2(new_n281), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n655), .A2(KEYINPUT15), .B1(new_n286), .B2(new_n288), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n299), .B1(new_n656), .B2(new_n298), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n296), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n296), .ZN(new_n660));
  NAND2_X1  g459(.A1(G229gat), .A2(G233gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT91), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n226), .B1(new_n297), .B2(new_n300), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT91), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n665), .A3(new_n660), .A4(new_n661), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT18), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n661), .B(KEYINPUT13), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n226), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n660), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n659), .A2(new_n662), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g474(.A(G113gat), .B(G141gat), .ZN(new_n676));
  INV_X1    g475(.A(G197gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT11), .B(G169gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT12), .Z(new_n681));
  NAND4_X1  g480(.A1(new_n663), .A2(new_n666), .A3(KEYINPUT92), .A4(new_n667), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n670), .A2(new_n675), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n675), .ZN(new_n684));
  INV_X1    g483(.A(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  AND4_X1   g486(.A1(new_n325), .A2(new_n634), .A3(new_n652), .A4(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n586), .A2(new_n587), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT100), .B(G1gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1324gat));
  NAND2_X1  g493(.A1(new_n688), .A2(new_n417), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G8gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT102), .Z(new_n697));
  XOR2_X1   g496(.A(KEYINPUT101), .B(KEYINPUT16), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G8gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n688), .A2(new_n417), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT42), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1325gat));
  NOR2_X1   g501(.A1(new_n542), .A2(new_n543), .ZN(new_n703));
  AOI21_X1  g502(.A(G15gat), .B1(new_n688), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n630), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n688), .B2(new_n706), .ZN(G1326gat));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n579), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NAND2_X1  g509(.A1(new_n634), .A2(new_n323), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n687), .A2(new_n322), .A3(new_n652), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n278), .A3(new_n691), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n625), .A2(new_n614), .B1(new_n631), .B2(new_n579), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n630), .A2(new_n716), .B1(new_n582), .B2(new_n598), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n717), .B2(new_n317), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n317), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n315), .A2(KEYINPUT104), .A3(new_n316), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n634), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n712), .B(KEYINPUT103), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n691), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1328gat));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n279), .A3(new_n417), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT46), .Z(new_n736));
  OAI21_X1  g535(.A(G36gat), .B1(new_n729), .B2(new_n583), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1329gat));
  NOR3_X1   g537(.A1(new_n729), .A2(new_n267), .A3(new_n630), .ZN(new_n739));
  AOI21_X1  g538(.A(G43gat), .B1(new_n713), .B2(new_n703), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g541(.A(new_n719), .B1(new_n634), .B2(new_n323), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT44), .B(new_n723), .C1(new_n599), .C2(new_n633), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n579), .B(new_n728), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n746), .A3(G50gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n746), .B1(new_n745), .B2(G50gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n713), .A2(new_n270), .A3(new_n579), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT48), .A4(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n726), .A2(KEYINPUT107), .A3(new_n579), .A4(new_n728), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(G50gat), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n757), .B2(new_n750), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT108), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n750), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT48), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762));
  INV_X1    g561(.A(new_n749), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n753), .A3(new_n750), .A4(new_n747), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n759), .A2(new_n765), .ZN(G1331gat));
  INV_X1    g565(.A(new_n687), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n325), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n651), .A3(new_n634), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n768), .A2(KEYINPUT109), .A3(new_n651), .A4(new_n634), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n691), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n205), .ZN(G1332gat));
  AND2_X1   g576(.A1(new_n771), .A2(new_n772), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT49), .B(G64gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n417), .A3(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n773), .A2(new_n583), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1333gat));
  INV_X1    g583(.A(new_n703), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n705), .A2(G71gat), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n786), .A2(G71gat), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n778), .A2(new_n579), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g591(.A1(new_n767), .A2(new_n322), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n711), .B2(new_n793), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n794), .A2(new_n691), .A3(new_n651), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n260), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n726), .A2(new_n322), .A3(new_n651), .A4(new_n767), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n691), .A2(G85gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT113), .ZN(G1336gat));
  AND2_X1   g600(.A1(new_n794), .A2(new_n795), .ZN(new_n802));
  INV_X1    g601(.A(G92gat), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n651), .A4(new_n417), .ZN(new_n804));
  INV_X1    g603(.A(new_n259), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n798), .B2(new_n583), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n798), .B2(new_n630), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n802), .A2(new_n651), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n785), .A2(G99gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(G1338gat));
  OAI21_X1  g611(.A(G106gat), .B1(new_n798), .B2(new_n596), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n596), .A2(G106gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT53), .ZN(G1339gat));
  AND4_X1   g615(.A1(new_n324), .A2(new_n318), .A3(new_n652), .A4(new_n767), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n682), .A2(new_n675), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n685), .B1(new_n668), .B2(new_n669), .ZN(new_n820));
  INV_X1    g619(.A(new_n680), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n660), .A2(new_n672), .A3(new_n671), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n664), .A2(new_n660), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n661), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n819), .A2(new_n820), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n643), .A2(new_n644), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n635), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n643), .A2(new_n636), .A3(new_n644), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n650), .B(new_n828), .C1(new_n830), .C2(new_n645), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n831), .A2(new_n832), .B1(new_n647), .B2(new_n650), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  INV_X1    g633(.A(new_n831), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(KEYINPUT55), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n832), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n825), .A2(new_n721), .A3(new_n722), .A4(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n821), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n683), .A2(new_n651), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n825), .A2(KEYINPUT115), .A3(new_n651), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n687), .A2(new_n838), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n840), .B1(new_n847), .B2(new_n723), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n818), .B1(new_n848), .B2(new_n252), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n580), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n691), .A2(new_n583), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n767), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n850), .A2(new_n417), .A3(new_n775), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n687), .A2(new_n437), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(G1340gat));
  OAI21_X1  g658(.A(G120gat), .B1(new_n852), .B2(new_n652), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n651), .B1(new_n435), .B2(new_n434), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n857), .B2(new_n861), .ZN(G1341gat));
  NAND2_X1  g661(.A1(new_n452), .A2(new_n448), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n852), .A2(new_n863), .A3(new_n322), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n854), .A2(new_n252), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n863), .ZN(G1342gat));
  OAI21_X1  g665(.A(G134gat), .B1(new_n852), .B2(new_n317), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n323), .A2(new_n583), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n850), .A2(G134gat), .A3(new_n775), .A4(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n870), .B2(new_n868), .ZN(new_n873));
  OAI221_X1 g672(.A(new_n867), .B1(new_n868), .B2(new_n870), .C1(new_n872), .C2(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n849), .A2(new_n875), .A3(new_n579), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n835), .B2(KEYINPUT55), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n831), .A2(KEYINPUT119), .A3(new_n832), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n683), .A2(new_n686), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n833), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n880), .A2(new_n881), .B1(new_n651), .B2(new_n825), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n839), .B1(new_n882), .B2(new_n323), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n817), .B1(new_n883), .B2(new_n322), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT57), .B1(new_n884), .B2(new_n596), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n851), .A2(new_n705), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT118), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n876), .A2(new_n885), .A3(new_n687), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n775), .A2(new_n705), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n849), .A2(new_n890), .A3(new_n583), .A4(new_n579), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n767), .A2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n891), .B2(new_n893), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n889), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(new_n891), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n892), .ZN(new_n900));
  AND4_X1   g699(.A1(KEYINPUT121), .A2(new_n889), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT58), .B1(new_n888), .B2(G141gat), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(new_n902), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n897), .B1(new_n901), .B2(new_n903), .ZN(G1344gat));
  AOI21_X1  g703(.A(new_n875), .B1(new_n849), .B2(new_n579), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n579), .A2(new_n875), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n882), .A2(new_n323), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n825), .A2(new_n323), .A3(new_n838), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n322), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n910), .B2(new_n818), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n906), .A2(new_n651), .A3(new_n887), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n899), .B2(new_n651), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n885), .A2(new_n887), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n915), .A3(new_n876), .ZN(new_n918));
  OAI221_X1 g717(.A(new_n914), .B1(G148gat), .B2(new_n916), .C1(new_n652), .C2(new_n918), .ZN(G1345gat));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n876), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(new_n426), .A3(new_n322), .ZN(new_n921));
  AOI21_X1  g720(.A(G155gat), .B1(new_n899), .B2(new_n252), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  NOR2_X1   g722(.A1(new_n424), .A2(new_n425), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n920), .B2(new_n723), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n869), .A2(new_n924), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n849), .A2(new_n890), .A3(new_n579), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n775), .A2(new_n417), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n850), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n767), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n691), .A2(new_n583), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n850), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n342), .A3(new_n687), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n936), .ZN(G1348gat));
  AOI21_X1  g736(.A(G176gat), .B1(new_n935), .B2(new_n651), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n652), .A2(new_n343), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n930), .B2(new_n939), .ZN(G1349gat));
  OAI21_X1  g739(.A(G183gat), .B1(new_n931), .B2(new_n322), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n252), .A3(new_n334), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n941), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1350gat));
  AOI21_X1  g745(.A(new_n333), .B1(new_n930), .B2(new_n323), .ZN(new_n947));
  XOR2_X1   g746(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  INV_X1    g750(.A(new_n935), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(G190gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n724), .ZN(new_n954));
  NOR4_X1   g753(.A1(new_n952), .A2(KEYINPUT123), .A3(G190gat), .A4(new_n723), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n949), .B(new_n950), .C1(new_n954), .C2(new_n955), .ZN(G1351gat));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n906), .A2(new_n957), .A3(new_n912), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n929), .A2(new_n705), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT125), .B1(new_n905), .B2(new_n911), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n767), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n849), .A2(new_n630), .A3(new_n579), .A4(new_n933), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n677), .A3(new_n687), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1352gat));
  XNOR2_X1  g765(.A(KEYINPUT126), .B(G204gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n967), .B1(new_n961), .B2(new_n652), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n963), .A2(new_n652), .ZN(new_n969));
  INV_X1    g768(.A(new_n967), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n972));
  NOR4_X1   g771(.A1(new_n963), .A2(KEYINPUT127), .A3(new_n652), .A4(new_n967), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n972), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n977), .B1(new_n969), .B2(new_n970), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n978), .B2(new_n973), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n968), .A2(new_n975), .A3(new_n979), .ZN(G1353gat));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n379), .A3(new_n252), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n906), .A2(new_n252), .A3(new_n912), .A4(new_n959), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(G218gat), .B1(new_n961), .B2(new_n317), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n964), .A2(new_n380), .A3(new_n724), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1355gat));
endmodule


