//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G58), .ZN(new_n205));
  INV_X1    g0005(.A(G232), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g0009(.A1(G107), .A2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n209), .B(new_n210), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n218), .B1(new_n217), .B2(new_n216), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(G50), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n224), .B(new_n227), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT65), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n228), .ZN(new_n254));
  NAND3_X1  g0054(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G226), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G223), .A2(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n269), .B(new_n270), .C1(G77), .C2(new_n265), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n264), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G200), .ZN(new_n274));
  INV_X1    g0074(.A(new_n273), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G190), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n228), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT67), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n257), .A2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G50), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  XOR2_X1   g0087(.A(KEYINPUT8), .B(G58), .Z(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT68), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n251), .A2(G20), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n289), .A2(new_n290), .B1(G150), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n229), .B1(new_n201), .B2(new_n212), .ZN(new_n293));
  XOR2_X1   g0093(.A(new_n293), .B(KEYINPUT69), .Z(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n287), .B1(new_n295), .B2(new_n279), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G50), .B2(new_n282), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n274), .B(new_n276), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n282), .A2(G50), .ZN(new_n300));
  AOI211_X1 g0100(.A(new_n300), .B(new_n287), .C1(new_n279), .C2(new_n295), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(KEYINPUT9), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n301), .A2(KEYINPUT9), .B1(G190), .B2(new_n275), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(new_n298), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n274), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n275), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n297), .B(new_n310), .C1(G169), .C2(new_n275), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(G58), .B(G68), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(G20), .B1(G159), .B2(new_n291), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT76), .B1(new_n315), .B2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(KEYINPUT76), .A3(G33), .ZN(new_n319));
  AOI21_X1  g0119(.A(G20), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(G68), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  OAI211_X1 g0123(.A(KEYINPUT16), .B(new_n314), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n321), .B1(new_n265), .B2(G20), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n315), .A2(G33), .ZN(new_n327));
  OAI211_X1 g0127(.A(KEYINPUT7), .B(new_n229), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT77), .B1(new_n329), .B2(G68), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT77), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  AOI211_X1 g0132(.A(new_n331), .B(new_n332), .C1(new_n325), .C2(new_n328), .ZN(new_n333));
  INV_X1    g0133(.A(new_n314), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n278), .B(new_n324), .C1(new_n335), .C2(KEYINPUT16), .ZN(new_n336));
  INV_X1    g0136(.A(new_n270), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n213), .A2(G1698), .ZN(new_n338));
  OR2_X1    g0138(.A1(G223), .A2(G1698), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n318), .A2(new_n338), .A3(new_n319), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n256), .A2(G232), .A3(new_n258), .ZN(new_n343));
  OR3_X1    g0143(.A1(new_n342), .A2(new_n343), .A3(new_n261), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(G200), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT8), .B(G58), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT68), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n257), .B2(G20), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n284), .B1(new_n283), .B2(new_n349), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n336), .A2(new_n346), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT17), .ZN(new_n353));
  NOR4_X1   g0153(.A1(new_n342), .A2(new_n343), .A3(new_n309), .A4(new_n261), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(G169), .B2(new_n344), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n336), .B2(new_n351), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT18), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT18), .ZN(new_n358));
  INV_X1    g0158(.A(new_n351), .ZN(new_n359));
  INV_X1    g0159(.A(new_n278), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n317), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n362), .B2(new_n229), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n321), .B(G20), .C1(new_n317), .C2(new_n361), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n331), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n329), .A2(KEYINPUT77), .A3(G68), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n314), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n360), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n359), .B1(new_n370), .B2(new_n324), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n358), .B1(new_n371), .B2(new_n355), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n256), .A2(new_n258), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n262), .B1(new_n374), .B2(new_n215), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT70), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G238), .A2(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n265), .B(new_n377), .C1(new_n206), .C2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n270), .C1(G107), .C2(new_n265), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  INV_X1    g0184(.A(new_n291), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n348), .A2(new_n385), .B1(new_n229), .B2(new_n214), .ZN(new_n386));
  XOR2_X1   g0186(.A(KEYINPUT15), .B(G87), .Z(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n290), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n384), .A2(new_n386), .B1(new_n388), .B2(KEYINPUT72), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n388), .A2(KEYINPUT72), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n384), .C2(new_n386), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n278), .B1(new_n214), .B2(new_n283), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n360), .A2(G77), .A3(new_n285), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n380), .B2(new_n345), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n353), .B(new_n373), .C1(new_n383), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n256), .A2(G238), .A3(new_n258), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G226), .A2(G1698), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n206), .B2(G1698), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(new_n265), .B1(G33), .B2(G97), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n399), .B(new_n262), .C1(new_n402), .C2(new_n337), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n398), .B1(new_n403), .B2(KEYINPUT13), .ZN(new_n404));
  INV_X1    g0204(.A(new_n403), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT74), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n408), .A3(KEYINPUT13), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n403), .B2(KEYINPUT13), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n404), .B(new_n407), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(G169), .C1(KEYINPUT75), .C2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n399), .A2(new_n262), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n406), .C1(new_n337), .C2(new_n402), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(G179), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n412), .A2(G169), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT75), .B(KEYINPUT14), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n414), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n290), .A2(G77), .B1(new_n291), .B2(G50), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n229), .B2(G68), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n279), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n424), .A2(KEYINPUT11), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n281), .A2(G20), .A3(new_n332), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT12), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(KEYINPUT11), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n360), .A2(G68), .A3(new_n285), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n425), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n416), .A2(G190), .A3(new_n417), .ZN(new_n432));
  AOI211_X1 g0232(.A(new_n430), .B(new_n432), .C1(new_n412), .C2(G200), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n381), .A2(new_n309), .ZN(new_n436));
  INV_X1    g0236(.A(G169), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n380), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n394), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n312), .A2(new_n397), .A3(new_n435), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n282), .A2(G97), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n325), .B2(new_n328), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n291), .A2(G77), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT6), .A2(G97), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G107), .ZN(new_n449));
  XNOR2_X1  g0249(.A(G97), .B(G107), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT6), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n447), .B1(new_n452), .B2(new_n229), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n446), .A2(KEYINPUT78), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n445), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT79), .B1(new_n455), .B2(new_n360), .ZN(new_n456));
  OAI21_X1  g0256(.A(G107), .B1(new_n363), .B2(new_n364), .ZN(new_n457));
  INV_X1    g0257(.A(new_n454), .ZN(new_n458));
  AND2_X1   g0258(.A1(G97), .A2(G107), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n451), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n444), .A2(KEYINPUT6), .A3(G97), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n463), .A2(G20), .B1(KEYINPUT78), .B2(new_n446), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n278), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n443), .B1(new_n456), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n257), .A2(G33), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n360), .A2(KEYINPUT67), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n277), .A2(KEYINPUT67), .A3(new_n228), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n282), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G97), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(G274), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n266), .A2(G244), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT76), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(KEYINPUT3), .B2(new_n251), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n319), .B(new_n481), .C1(new_n483), .C2(new_n326), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n480), .A2(new_n485), .B1(new_n208), .B2(new_n266), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n265), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n479), .B1(new_n490), .B2(new_n270), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n475), .A2(new_n477), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n256), .A3(G257), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(G190), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n493), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n468), .A2(new_n474), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n443), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n465), .A2(new_n466), .A3(new_n278), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n466), .B1(new_n465), .B2(new_n278), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n474), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n437), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n491), .A2(new_n309), .A3(new_n493), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n266), .A2(G264), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n220), .A2(new_n266), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n318), .A2(new_n319), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n362), .A2(G303), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n337), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n492), .A2(new_n256), .A3(G270), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n511), .A2(new_n479), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n257), .A2(new_n514), .A3(G13), .A4(G20), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n360), .A2(new_n282), .A3(G116), .A4(new_n469), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n277), .A2(new_n228), .B1(G20), .B2(new_n514), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n487), .B(new_n229), .C1(G33), .C2(new_n219), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n519), .A2(KEYINPUT20), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT20), .B1(new_n519), .B2(new_n520), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n517), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n513), .A2(G179), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n513), .A2(G190), .ZN(new_n525));
  INV_X1    g0325(.A(new_n523), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(new_n382), .C2(new_n513), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n513), .A2(new_n437), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n523), .ZN(new_n530));
  NOR4_X1   g0330(.A1(new_n513), .A2(new_n526), .A3(KEYINPUT21), .A4(new_n437), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n524), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n215), .A2(G1698), .ZN(new_n533));
  OR2_X1    g0333(.A1(G238), .A2(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n318), .A2(new_n319), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n270), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n477), .A2(G274), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n256), .B(G250), .C1(G1), .C2(new_n476), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G200), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(G190), .A3(new_n542), .A4(new_n543), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n318), .A2(new_n319), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n229), .A3(G68), .ZN(new_n548));
  NOR3_X1   g0348(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(G33), .B2(G97), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT19), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OR3_X1    g0351(.A1(new_n251), .A2(new_n219), .A3(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(G20), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n360), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n472), .A2(new_n207), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n387), .A2(new_n282), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n545), .A2(new_n546), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n544), .A2(G169), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n541), .A2(G179), .A3(new_n542), .A4(new_n543), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n554), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n473), .A2(new_n387), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n532), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n220), .A2(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n208), .A2(new_n266), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n318), .A2(new_n319), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G294), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n337), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n492), .A2(new_n256), .A3(G264), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(new_n479), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT84), .B1(new_n571), .B2(new_n437), .ZN(new_n572));
  INV_X1    g0372(.A(new_n570), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n567), .A2(new_n568), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n478), .C1(new_n574), .C2(new_n337), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(G169), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(G179), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n207), .A2(G20), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n317), .A3(new_n361), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n229), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n444), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n581), .A2(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n318), .A2(KEYINPUT22), .A3(new_n319), .A4(new_n580), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n290), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT83), .A4(new_n588), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(KEYINPUT24), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT24), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n278), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n281), .A2(G20), .A3(new_n444), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n473), .B2(G107), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n579), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n571), .A2(G190), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n575), .A2(G200), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n596), .A2(new_n599), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT80), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n497), .A2(new_n504), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n506), .A2(new_n564), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n442), .A2(new_n609), .ZN(G372));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n371), .A2(new_n358), .A3(new_n355), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n336), .A2(new_n351), .ZN(new_n613));
  INV_X1    g0413(.A(new_n355), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT18), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n357), .A2(new_n372), .A3(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n431), .B1(new_n433), .B2(new_n439), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n353), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n308), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n311), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n561), .A2(new_n562), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n559), .A2(new_n626), .A3(new_n560), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n559), .B2(new_n560), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n504), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n559), .A2(new_n560), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n625), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n546), .A2(new_n557), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n545), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n604), .ZN(new_n641));
  INV_X1    g0441(.A(new_n524), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n511), .A2(new_n512), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n478), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(G169), .A3(new_n523), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT21), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n529), .A2(new_n528), .A3(new_n523), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n641), .B1(new_n648), .B2(new_n601), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n634), .B1(new_n649), .B2(new_n497), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT86), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n545), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n544), .A2(KEYINPUT86), .A3(G200), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n637), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n629), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n633), .B(new_n640), .C1(new_n650), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n624), .B1(new_n442), .B2(new_n658), .ZN(G369));
  OAI21_X1  g0459(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n280), .A2(G20), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n257), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n526), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n532), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT89), .B(G330), .Z(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n668), .B1(new_n596), .B2(new_n599), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n605), .A2(new_n675), .B1(new_n601), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n605), .A2(new_n648), .A3(new_n667), .ZN(new_n678));
  INV_X1    g0478(.A(new_n601), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n668), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n225), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G1), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n549), .A2(new_n514), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n232), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n633), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n559), .A2(new_n626), .A3(new_n560), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n653), .A2(new_n654), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n694), .A2(new_n625), .B1(new_n695), .B2(new_n637), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n505), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n497), .A2(new_n504), .A3(KEYINPUT93), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n696), .A2(new_n649), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n639), .A2(new_n651), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n629), .A2(KEYINPUT26), .A3(new_n634), .A4(new_n655), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n630), .A2(KEYINPUT92), .A3(new_n632), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n691), .A2(new_n700), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n689), .B1(new_n705), .B2(new_n668), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n657), .A2(new_n668), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT91), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT91), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n657), .A2(new_n709), .A3(new_n668), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n706), .B1(new_n711), .B2(new_n689), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n491), .A2(new_n571), .A3(new_n643), .A4(new_n493), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n560), .ZN(new_n715));
  NOR2_X1   g0515(.A1(KEYINPUT90), .A2(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n571), .A2(G179), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n544), .A2(new_n719), .A3(new_n495), .A4(new_n644), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n716), .B1(new_n713), .B2(new_n560), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n667), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n725), .A3(new_n667), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n609), .B2(new_n667), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n672), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT94), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n688), .B1(new_n731), .B2(G1), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT95), .ZN(G364));
  NAND2_X1  g0533(.A1(new_n661), .A2(G45), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n684), .A2(G1), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT96), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n229), .A2(new_n345), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n382), .A2(G179), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G87), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n309), .A2(new_n382), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n229), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n737), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n741), .B1(new_n744), .B2(new_n332), .C1(new_n212), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n738), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n265), .B1(new_n747), .B2(new_n444), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n219), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n746), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n743), .A2(new_n749), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n309), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n737), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n743), .A2(new_n759), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n205), .B1(new_n761), .B2(new_n214), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT98), .Z(new_n763));
  NAND3_X1  g0563(.A1(new_n754), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT99), .Z(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n747), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n362), .B1(new_n739), .B2(new_n768), .C1(new_n769), .C2(new_n760), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(G294), .B2(new_n751), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n745), .A2(new_n772), .B1(new_n761), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n755), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G329), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n744), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n771), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n765), .B1(new_n767), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n228), .B1(G20), .B2(new_n437), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n736), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n265), .A2(G355), .A3(new_n225), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n547), .A2(new_n682), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G45), .B2(new_n232), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n245), .A2(new_n476), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n786), .B1(G116), .B2(new_n225), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n229), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  INV_X1    g0593(.A(new_n784), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n785), .B(new_n796), .C1(new_n671), .C2(new_n793), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n671), .A2(new_n672), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n673), .A3(new_n735), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(G396));
  NOR2_X1   g0600(.A1(new_n439), .A2(new_n667), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n396), .A2(new_n383), .B1(new_n395), .B2(new_n668), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n439), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n657), .A2(new_n668), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n711), .B2(new_n803), .ZN(new_n805));
  INV_X1    g0605(.A(new_n672), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n636), .A2(new_n638), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(new_n605), .A3(new_n532), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n808), .A2(new_n506), .A3(new_n608), .A4(new_n668), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(new_n809), .B2(new_n727), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n805), .B(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(new_n735), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n784), .A2(new_n791), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G77), .ZN(new_n815));
  INV_X1    g0615(.A(new_n736), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n747), .A2(new_n207), .ZN(new_n817));
  INV_X1    g0617(.A(new_n760), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G294), .B2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n819), .B1(new_n514), .B2(new_n761), .C1(new_n768), .C2(new_n745), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n739), .A2(new_n444), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n362), .B1(new_n755), .B2(new_n773), .C1(new_n766), .C2(new_n744), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n820), .A2(new_n753), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G143), .A2(new_n818), .B1(new_n777), .B2(G150), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n825), .B2(new_n745), .C1(new_n756), .C2(new_n761), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT34), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n547), .B1(new_n205), .B2(new_n752), .ZN(new_n828));
  INV_X1    g0628(.A(new_n747), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G68), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n212), .B2(new_n739), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n827), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n775), .A2(G132), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n823), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n816), .B1(new_n834), .B2(new_n794), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n802), .A2(new_n439), .ZN(new_n836));
  INV_X1    g0636(.A(new_n801), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n815), .B(new_n835), .C1(new_n791), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n812), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  OAI211_X1 g0641(.A(G116), .B(new_n230), .C1(new_n463), .C2(KEYINPUT35), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT100), .Z(new_n843));
  INV_X1    g0643(.A(KEYINPUT35), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n452), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT36), .ZN(new_n846));
  OAI21_X1  g0646(.A(G77), .B1(new_n205), .B2(new_n332), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n232), .A2(new_n847), .B1(G50), .B2(new_n332), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(G1), .A3(new_n280), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT101), .Z(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT104), .B1(new_n712), .B2(new_n442), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n604), .B(new_n497), .C1(new_n679), .C2(new_n660), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n504), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n651), .A3(new_n696), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n630), .A2(new_n632), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n856));
  AOI211_X1 g0656(.A(KEYINPUT91), .B(new_n667), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n709), .B1(new_n657), .B2(new_n668), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n689), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n706), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT104), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n441), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n623), .B1(new_n852), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n314), .B1(new_n322), .B2(new_n323), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n369), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n279), .A3(new_n324), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n351), .ZN(new_n869));
  INV_X1    g0669(.A(new_n665), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n869), .B1(new_n614), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n865), .B1(new_n871), .B2(new_n352), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n352), .B1(new_n371), .B2(new_n355), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT102), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n371), .B2(new_n665), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n613), .A2(KEYINPUT102), .A3(new_n870), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(new_n865), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n336), .A2(new_n347), .A3(new_n351), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n356), .B1(new_n882), .B2(new_n346), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n883), .A3(new_n874), .A4(new_n865), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n873), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n869), .A2(new_n870), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n353), .B2(new_n373), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n881), .A2(new_n883), .A3(new_n865), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n872), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n891), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n804), .A2(new_n837), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n430), .A2(new_n667), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n431), .A2(new_n434), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n430), .B(new_n667), .C1(new_n421), .C2(new_n433), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n880), .A2(new_n885), .B1(new_n865), .B2(new_n879), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n881), .B1(new_n618), .B2(new_n353), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n894), .A2(new_n891), .A3(new_n888), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n431), .A2(new_n667), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n890), .A2(new_n895), .A3(KEYINPUT39), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n619), .A2(new_n665), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n864), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n728), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n838), .B1(new_n899), .B2(new_n900), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n809), .A2(KEYINPUT105), .A3(new_n727), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n896), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n865), .B1(new_n881), .B2(new_n883), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n893), .B2(new_n884), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n891), .B1(new_n926), .B2(new_n906), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n890), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n809), .A2(KEYINPUT105), .A3(new_n727), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT105), .B1(new_n809), .B2(new_n727), .ZN(new_n930));
  INV_X1    g0730(.A(new_n900), .ZN(new_n931));
  INV_X1    g0731(.A(new_n898), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n433), .B(new_n932), .C1(new_n421), .C2(new_n430), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n803), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n928), .A2(KEYINPUT40), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n920), .A2(new_n922), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n442), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n672), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n917), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n661), .A2(new_n257), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n851), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OAI21_X1  g0744(.A(new_n265), .B1(new_n739), .B2(new_n205), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G77), .A2(new_n829), .B1(new_n775), .B2(G137), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n756), .B2(new_n744), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT111), .ZN(new_n948));
  INV_X1    g0748(.A(new_n745), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n949), .A2(G143), .B1(new_n751), .B2(G68), .ZN(new_n950));
  INV_X1    g0750(.A(G150), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n760), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n945), .B(new_n947), .C1(new_n948), .C2(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n948), .B2(new_n952), .C1(new_n212), .C2(new_n761), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n755), .A2(new_n778), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n829), .A2(G97), .ZN(new_n956));
  INV_X1    g0756(.A(G294), .ZN(new_n957));
  XOR2_X1   g0757(.A(KEYINPUT110), .B(G311), .Z(new_n958));
  OAI221_X1 g0758(.A(new_n956), .B1(new_n957), .B2(new_n744), .C1(new_n745), .C2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n761), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(G283), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n739), .A2(new_n514), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n962), .A2(KEYINPUT46), .B1(new_n752), .B2(new_n444), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT46), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n547), .B1(G303), .B2(new_n818), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n954), .B1(new_n955), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n736), .B1(new_n969), .B2(new_n784), .ZN(new_n970));
  INV_X1    g0770(.A(new_n387), .ZN(new_n971));
  INV_X1    g0771(.A(new_n787), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n795), .B1(new_n225), .B2(new_n971), .C1(new_n972), .C2(new_n241), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n696), .B1(new_n557), .B2(new_n668), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n557), .A2(new_n668), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n633), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n970), .B(new_n973), .C1(new_n976), .C2(new_n793), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n734), .A2(G1), .ZN(new_n978));
  INV_X1    g0778(.A(new_n677), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n501), .A2(new_n667), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n698), .A2(new_n699), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n504), .A2(new_n668), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT107), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(KEYINPUT107), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n680), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n987), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n985), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(KEYINPUT45), .A3(new_n680), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n992), .B2(new_n680), .ZN(new_n997));
  INV_X1    g0797(.A(new_n680), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n991), .A2(new_n998), .A3(new_n985), .A4(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n979), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n990), .A2(new_n993), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1002), .A2(new_n677), .A3(new_n999), .A4(new_n997), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n678), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n648), .A2(new_n667), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n676), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n673), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n731), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n683), .B(KEYINPUT41), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n978), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT42), .B1(new_n992), .B2(new_n678), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT42), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1013), .B(new_n1005), .C1(new_n991), .C2(new_n985), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT106), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT43), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n976), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT108), .B1(new_n986), .B2(new_n987), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT108), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n991), .A2(new_n1022), .A3(new_n985), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1023), .A3(new_n679), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1024), .A2(new_n504), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1016), .B(new_n1020), .C1(new_n1025), .C2(new_n667), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1020), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n667), .B1(new_n1024), .B2(new_n504), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(new_n1015), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n979), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1026), .A2(new_n1030), .A3(new_n979), .A4(new_n1032), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n977), .B1(new_n1011), .B2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n1008), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n747), .A2(new_n514), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n547), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G322), .A2(new_n949), .B1(new_n960), .B2(G303), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n778), .B2(new_n760), .C1(new_n744), .C2(new_n958), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT48), .Z(new_n1043));
  AOI22_X1  g0843(.A1(new_n740), .A2(G294), .B1(new_n751), .B2(G283), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1040), .B1(new_n772), .B2(new_n755), .C1(new_n1047), .C2(KEYINPUT49), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1039), .B(new_n1048), .C1(KEYINPUT49), .C2(new_n1047), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n740), .A2(G77), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n775), .A2(G150), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1050), .A2(new_n956), .A3(new_n547), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n752), .A2(new_n971), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n745), .A2(new_n756), .B1(new_n760), .B2(new_n212), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1054), .B(new_n1057), .C1(new_n349), .C2(new_n744), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1053), .B(new_n1058), .C1(G68), .C2(new_n960), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n784), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n676), .A2(new_n793), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n288), .A2(new_n212), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n686), .B1(new_n1062), .B2(KEYINPUT50), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(G68), .A2(G77), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n476), .A4(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n787), .B(new_n1066), .C1(new_n238), .C2(new_n476), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n686), .A2(new_n225), .A3(new_n265), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G107), .C2(new_n225), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT113), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n736), .B(new_n1061), .C1(new_n795), .C2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n978), .A2(new_n1038), .B1(new_n1060), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n683), .B1(new_n731), .B2(new_n1038), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT94), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n730), .B(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n1008), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1072), .B1(new_n1073), .B2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n731), .A2(new_n1038), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n684), .B1(new_n1078), .B2(new_n1004), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n731), .A2(new_n1003), .A3(new_n1001), .A4(new_n1038), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1001), .A2(new_n978), .A3(new_n1003), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n795), .B1(new_n219), .B2(new_n225), .C1(new_n972), .C2(new_n248), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n817), .B(new_n1040), .C1(G143), .C2(new_n775), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n745), .A2(new_n951), .B1(new_n760), .B2(new_n756), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n739), .A2(new_n332), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n744), .A2(new_n212), .B1(new_n761), .B2(new_n348), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G77), .C2(new_n751), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n745), .A2(new_n778), .B1(new_n760), .B2(new_n773), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n444), .B2(new_n747), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n744), .A2(new_n768), .B1(new_n761), .B2(new_n957), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G322), .B2(new_n775), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n751), .A2(G116), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n740), .A2(G283), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1095), .A2(new_n362), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1090), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n736), .B1(new_n1099), .B2(new_n784), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1083), .B(new_n1100), .C1(new_n1032), .C2(new_n793), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1082), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1081), .A2(new_n1103), .ZN(G390));
  NAND4_X1  g0904(.A1(new_n920), .A2(G330), .A3(new_n803), .A4(new_n922), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n901), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n911), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n910), .A2(new_n912), .B1(new_n1109), .B2(new_n902), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n928), .A2(new_n1109), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n705), .A2(new_n668), .A3(new_n836), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n1112), .B2(new_n837), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1108), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n902), .A2(new_n1109), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n912), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT39), .B1(new_n890), .B2(new_n927), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1112), .A2(new_n837), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1109), .B(new_n928), .C1(new_n1120), .C2(new_n1106), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n810), .A2(new_n803), .A3(new_n901), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT116), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT116), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n810), .A2(new_n1124), .A3(new_n803), .A4(new_n901), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1119), .A2(new_n1121), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n939), .A2(G330), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n862), .B1(new_n861), .B2(new_n441), .ZN(new_n1130));
  AOI211_X1 g0930(.A(KEYINPUT104), .B(new_n442), .C1(new_n859), .C2(new_n860), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n624), .B(new_n1129), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1126), .A2(new_n1120), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1106), .B1(new_n729), .B2(new_n838), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n897), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT117), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(KEYINPUT117), .A3(new_n897), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1115), .B(new_n1128), .C1(new_n1132), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1115), .A2(new_n1128), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1126), .A2(new_n1120), .A3(new_n1133), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1140), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT117), .B1(new_n1136), .B2(new_n897), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n864), .A3(new_n1129), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1148), .A3(new_n683), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n978), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1115), .B2(new_n1128), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT120), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n289), .A2(new_n814), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n777), .A2(G107), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n741), .A2(new_n1154), .A3(new_n830), .A4(new_n362), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G116), .A2(new_n818), .B1(new_n960), .B2(G97), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n766), .B2(new_n745), .C1(new_n957), .C2(new_n755), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G77), .C2(new_n751), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n362), .B1(new_n829), .B2(G50), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT119), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT118), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1160), .B1(new_n1163), .B2(new_n761), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G128), .A2(new_n949), .B1(new_n777), .B2(G137), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n755), .C1(KEYINPUT119), .C2(new_n1159), .ZN(new_n1167));
  INV_X1    g0967(.A(G132), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n760), .A2(new_n1168), .ZN(new_n1169));
  OR3_X1    g0969(.A1(new_n739), .A2(KEYINPUT53), .A3(new_n951), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT53), .B1(new_n739), .B2(new_n951), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n756), .C2(new_n752), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1164), .A2(new_n1167), .A3(new_n1169), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n784), .B1(new_n1158), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n816), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n910), .A2(new_n912), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1153), .B(new_n1175), .C1(new_n1176), .C2(new_n791), .ZN(new_n1177));
  OR3_X1    g0977(.A1(new_n1151), .A2(new_n1152), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1152), .B1(new_n1151), .B2(new_n1177), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1149), .A2(new_n1178), .A3(new_n1179), .ZN(G378));
  AOI21_X1  g0980(.A(new_n923), .B1(new_n890), .B2(new_n895), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n936), .B(G330), .C1(new_n1181), .C2(KEYINPUT40), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n312), .A2(KEYINPUT55), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT55), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n308), .B2(new_n311), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n297), .A2(new_n870), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT56), .Z(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1183), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1182), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n924), .A2(G330), .A3(new_n936), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n916), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT122), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1192), .A2(new_n915), .A3(new_n1194), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1132), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1110), .A2(new_n1114), .A3(new_n1126), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1107), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1200), .B1(new_n1203), .B2(new_n1141), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n915), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT122), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1199), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT57), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n684), .B1(new_n1210), .B2(new_n1204), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1199), .A2(new_n978), .A3(new_n1206), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G128), .A2(new_n818), .B1(new_n777), .B2(G132), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1166), .B2(new_n745), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G150), .B2(new_n751), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n825), .B2(new_n761), .C1(new_n739), .C2(new_n1163), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT59), .Z(new_n1218));
  AOI21_X1  g1018(.A(G41), .B1(new_n775), .B2(G124), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G33), .B1(new_n829), .B2(G159), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1040), .A2(new_n252), .A3(new_n1050), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT121), .Z(new_n1223));
  OAI22_X1  g1023(.A1(new_n971), .A2(new_n761), .B1(new_n766), .B2(new_n755), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G97), .B2(new_n777), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n205), .B2(new_n747), .C1(new_n444), .C2(new_n760), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n752), .A2(new_n332), .B1(new_n745), .B2(new_n514), .ZN(new_n1227));
  OR3_X1    g1027(.A1(new_n1223), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT58), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G41), .B1(new_n547), .B2(G33), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1221), .B(new_n1229), .C1(G50), .C2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n735), .B1(new_n1231), .B2(new_n784), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n791), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1232), .B1(G50), .B2(new_n814), .C1(new_n1191), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1213), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1212), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1106), .A2(new_n791), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n813), .A2(new_n332), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n362), .B1(new_n747), .B2(new_n214), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1240), .B(new_n1055), .C1(G303), .C2(new_n775), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n745), .A2(new_n957), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n760), .A2(new_n766), .B1(new_n761), .B2(new_n444), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G97), .C2(new_n740), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1241), .B(new_n1244), .C1(new_n514), .C2(new_n744), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n761), .A2(new_n951), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1040), .B1(G159), .B2(new_n740), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n829), .A2(G58), .B1(new_n751), .B2(G50), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1162), .A2(new_n777), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n745), .A2(new_n1168), .B1(new_n760), .B2(new_n825), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G128), .B2(new_n775), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1246), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n736), .B1(new_n1253), .B2(new_n784), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1238), .A2(new_n1239), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1141), .B2(new_n1150), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1010), .B1(new_n1200), .B2(new_n1147), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1132), .A2(new_n1141), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(G381));
  INV_X1    g1060(.A(G396), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1072), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(G384), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT123), .ZN(new_n1264));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1212), .A2(new_n1265), .A3(new_n1236), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1102), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1267), .B(new_n977), .C1(new_n1011), .C2(new_n1036), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G381), .A2(new_n1264), .A3(new_n1266), .A4(new_n1268), .ZN(G407));
  INV_X1    g1069(.A(G213), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1266), .A2(new_n1270), .A3(G343), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(G407), .A2(new_n1272), .A3(G213), .A4(new_n1273), .ZN(G409));
  AOI21_X1  g1074(.A(new_n1265), .B1(new_n1212), .B2(new_n1236), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1199), .A2(new_n1204), .A3(new_n1010), .A4(new_n1206), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1192), .A2(new_n915), .A3(new_n1194), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n978), .B1(new_n1277), .B2(new_n1205), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1149), .A2(new_n1178), .A3(new_n1179), .A4(new_n1234), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1279), .A2(new_n1280), .B1(new_n1270), .B2(G343), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT126), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT60), .B1(new_n1132), .B2(new_n1141), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1283), .A2(new_n1259), .A3(new_n684), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1132), .A2(new_n1141), .A3(KEYINPUT60), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1132), .A2(new_n1141), .A3(KEYINPUT125), .A4(KEYINPUT60), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1257), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n840), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(G384), .A3(new_n1257), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1270), .A2(G343), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1290), .B2(new_n1257), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n840), .B(new_n1256), .C1(new_n1284), .C2(new_n1289), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1295), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1205), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1132), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n683), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1208), .B2(new_n1207), .ZN(new_n1305));
  OAI21_X1  g1105(.A(G378), .B1(new_n1305), .B2(new_n1235), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1280), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1294), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1306), .A2(new_n1307), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1282), .A2(new_n1301), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1306), .A2(new_n1314), .A3(new_n1310), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1306), .A2(new_n1314), .A3(new_n1310), .A4(KEYINPUT63), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1312), .A2(new_n1313), .A3(new_n1317), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G387), .A2(G390), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G393), .A2(G396), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1262), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1320), .A2(new_n1268), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1320), .B2(new_n1268), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1315), .A2(new_n1326), .ZN(new_n1327));
  OR2_X1    g1127(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1306), .A2(new_n1314), .A3(new_n1310), .A4(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1325), .B1(new_n1331), .B2(new_n1301), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1319), .A2(new_n1325), .B1(new_n1330), .B2(new_n1332), .ZN(G405));
  INV_X1    g1133(.A(new_n1266), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1314), .B1(new_n1334), .B2(new_n1275), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1306), .B(new_n1266), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1337), .B(new_n1325), .ZN(G402));
endmodule


