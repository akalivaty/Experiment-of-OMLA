//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OR3_X1    g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n210), .B(new_n213), .C1(KEYINPUT15), .C2(new_n207), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(KEYINPUT91), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n211), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n212), .A2(KEYINPUT91), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT15), .A3(new_n207), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G1gat), .B2(new_n222), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT93), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n214), .A2(new_n220), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n227), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT13), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n232), .A2(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n227), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n231), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n235), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT18), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n206), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n237), .B(KEYINPUT94), .ZN(new_n248));
  INV_X1    g047(.A(new_n206), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n245), .B(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G211gat), .B(G218gat), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  XOR2_X1   g055(.A(G197gat), .B(G204gat), .Z(new_n257));
  AOI21_X1  g056(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n256), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT79), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n261), .A2(new_n262), .B1(G155gat), .B2(G162gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n264));
  INV_X1    g063(.A(G141gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G148gat), .ZN(new_n266));
  INV_X1    g065(.A(G148gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G141gat), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n263), .A2(new_n264), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT78), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G155gat), .A3(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G155gat), .ZN(new_n275));
  INV_X1    g074(.A(G162gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT80), .B1(new_n269), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n270), .B1(KEYINPUT79), .B2(KEYINPUT2), .ZN(new_n280));
  INV_X1    g079(.A(new_n264), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n267), .A2(G141gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n265), .A2(G148gat), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n271), .A2(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT81), .B1(new_n265), .B2(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(new_n267), .A3(G141gat), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT82), .A4(new_n266), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n266), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n262), .A2(new_n275), .A3(new_n276), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n292), .A2(new_n293), .B1(new_n270), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n287), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n260), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n259), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n254), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n259), .A2(KEYINPUT86), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(new_n304), .A3(new_n255), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n299), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n297), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n293), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n270), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n291), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT83), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n279), .A2(new_n287), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT83), .A3(new_n313), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n256), .B(new_n303), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n297), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n300), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n318), .B1(new_n326), .B2(new_n302), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G22gat), .ZN(new_n328));
  INV_X1    g127(.A(G22gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n318), .B(new_n329), .C1(new_n326), .C2(new_n302), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G78gat), .B(G106gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G50gat), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n335), .B(new_n336), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n328), .A2(new_n330), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G113gat), .ZN(new_n343));
  INV_X1    g142(.A(G120gat), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT1), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G134gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(G127gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G134gat), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n352));
  OAI21_X1  g151(.A(G120gat), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n345), .B1(new_n343), .B2(new_n344), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n349), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n350), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n320), .A2(new_n322), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n313), .B(new_n356), .C1(new_n314), .C2(new_n315), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT39), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n320), .A2(KEYINPUT3), .A3(new_n322), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n356), .B1(new_n296), .B2(new_n297), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n321), .A2(KEYINPUT4), .A3(new_n313), .A4(new_n356), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n361), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT0), .ZN(new_n374));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT39), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n372), .A2(KEYINPUT40), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT40), .B1(new_n372), .B2(new_n379), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n368), .A2(new_n361), .A3(new_n369), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n366), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n362), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n366), .A3(new_n386), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n380), .A2(new_n381), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G226gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n395));
  INV_X1    g194(.A(G169gat), .ZN(new_n396));
  INV_X1    g195(.A(G176gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT23), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(KEYINPUT23), .ZN(new_n403));
  NOR2_X1   g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT24), .ZN(new_n405));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n395), .B1(new_n400), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT69), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT67), .B(KEYINPUT24), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n406), .B1(new_n412), .B2(new_n404), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n408), .B(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT25), .B1(new_n402), .B2(KEYINPUT23), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n398), .A2(KEYINPUT66), .A3(new_n401), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT66), .B1(new_n398), .B2(new_n401), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n413), .A2(new_n411), .A3(new_n415), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n410), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G183gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT27), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT27), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G183gat), .ZN(new_n428));
  INV_X1    g227(.A(G190gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT28), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT27), .B(G183gat), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT28), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n429), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n434), .A3(new_n406), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT70), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n436), .A2(new_n437), .A3(new_n401), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n436), .B2(new_n401), .ZN(new_n439));
  NOR3_X1   g238(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT75), .B(new_n394), .C1(new_n424), .C2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT75), .ZN(new_n444));
  INV_X1    g243(.A(new_n406), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n405), .A2(KEYINPUT67), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT24), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n404), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n408), .B(KEYINPUT68), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT69), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n398), .A2(new_n401), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT66), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n398), .A2(KEYINPUT66), .A3(new_n401), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n417), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(new_n458), .A3(new_n423), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n400), .A2(new_n409), .ZN(new_n460));
  INV_X1    g259(.A(new_n395), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n442), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n394), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n444), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n443), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n463), .B2(KEYINPUT29), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n260), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n459), .A2(new_n462), .ZN(new_n469));
  INV_X1    g268(.A(new_n442), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n394), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n467), .A3(new_n260), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(G64gat), .B(G92gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT76), .B1(new_n468), .B2(new_n474), .ZN(new_n482));
  INV_X1    g281(.A(new_n478), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n299), .B1(new_n424), .B2(new_n442), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n443), .A2(new_n465), .B1(new_n485), .B2(new_n464), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n484), .B(new_n473), .C1(new_n486), .C2(new_n260), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n342), .B1(new_n391), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n382), .B1(new_n364), .B2(new_n365), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n361), .B1(new_n358), .B2(new_n359), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n495), .A2(new_n386), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n389), .A2(new_n376), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n499), .B2(new_n390), .ZN(new_n500));
  INV_X1    g299(.A(new_n389), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n377), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n377), .B1(new_n495), .B2(new_n386), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT6), .B1(new_n503), .B2(new_n388), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(new_n473), .C1(new_n486), .C2(new_n260), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n472), .A2(new_n467), .A3(new_n324), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT37), .B(new_n509), .C1(new_n486), .C2(new_n324), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT38), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(new_n483), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT6), .B(new_n377), .C1(new_n497), .C2(new_n501), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n479), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n492), .B1(new_n506), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n512), .A2(new_n513), .A3(new_n479), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n516), .A2(KEYINPUT89), .A3(new_n500), .A4(new_n505), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n482), .A2(KEYINPUT37), .A3(new_n487), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n508), .A2(new_n483), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n491), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n471), .A2(new_n356), .ZN(new_n525));
  NAND2_X1  g324(.A1(G227gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n463), .A2(new_n357), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT32), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G15gat), .B(G43gat), .Z(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n529), .B(KEYINPUT32), .C1(new_n531), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n528), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(new_n526), .ZN(new_n543));
  AOI211_X1 g342(.A(new_n527), .B(new_n540), .C1(new_n525), .C2(new_n528), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n536), .B(new_n538), .C1(new_n544), .C2(new_n543), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT36), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n546), .A3(new_n547), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n539), .A2(KEYINPUT73), .A3(new_n545), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n552), .B2(KEYINPUT36), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n488), .A2(KEYINPUT77), .A3(new_n489), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n513), .B1(new_n499), .B2(new_n390), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n481), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT77), .B1(new_n488), .B2(new_n489), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n342), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n524), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n546), .A2(new_n547), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n342), .A2(new_n562), .A3(KEYINPUT35), .ZN(new_n563));
  INV_X1    g362(.A(new_n490), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n500), .A2(new_n505), .A3(new_n513), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n557), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(new_n555), .A3(new_n481), .A4(new_n554), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n341), .A2(new_n550), .A3(new_n551), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT35), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n253), .B1(new_n560), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G230gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n393), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(G85gat), .A3(G92gat), .ZN(new_n577));
  INV_X1    g376(.A(G85gat), .ZN(new_n578));
  INV_X1    g377(.A(G92gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n581), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G99gat), .B(G106gat), .Z(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n588));
  XNOR2_X1  g387(.A(G57gat), .B(G64gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n587), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR3_X1    g395(.A1(new_n587), .A2(new_n595), .A3(new_n593), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n574), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n594), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n574), .ZN(new_n600));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  OR2_X1    g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n574), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n241), .A2(new_n587), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(new_n240), .ZN(new_n611));
  INV_X1    g410(.A(new_n587), .ZN(new_n612));
  AND2_X1   g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n612), .A2(new_n221), .B1(KEYINPUT41), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  OR3_X1    g415(.A1(new_n615), .A2(KEYINPUT101), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT101), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT98), .ZN(new_n620));
  XOR2_X1   g419(.A(G134gat), .B(G162gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n616), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n617), .A2(new_n618), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(KEYINPUT99), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n615), .A2(new_n616), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n227), .B1(new_n630), .B2(new_n593), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n593), .A2(new_n630), .ZN(new_n633));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n632), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n636), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n572), .A2(new_n609), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n555), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n564), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n226), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n226), .B2(new_n651), .ZN(new_n655));
  MUX2_X1   g454(.A(new_n654), .B(new_n655), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n648), .B2(new_n553), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n562), .A2(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n648), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n648), .A2(new_n341), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT103), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n560), .A2(new_n571), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n609), .A2(new_n646), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n253), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n629), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n555), .A2(G29gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n665), .B2(new_n629), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n629), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n624), .A2(KEYINPUT106), .A3(new_n628), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n558), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n568), .A2(KEYINPUT105), .A3(new_n342), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n524), .A2(new_n553), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n684), .B2(new_n571), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n667), .B1(new_n676), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT107), .B(new_n667), .C1(new_n676), .C2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n555), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n664), .B1(new_n674), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n672), .B(KEYINPUT45), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(KEYINPUT108), .A3(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1328gat));
  OAI21_X1  g495(.A(G36gat), .B1(new_n690), .B2(new_n564), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n668), .A2(G36gat), .A3(new_n564), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(G1329gat));
  OAI21_X1  g499(.A(G43gat), .B1(new_n686), .B2(new_n553), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n668), .A2(G43gat), .A3(new_n562), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n553), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n688), .A2(new_n706), .A3(new_n689), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n707), .A2(KEYINPUT109), .A3(G43gat), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT109), .B1(new_n707), .B2(G43gat), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n708), .A2(new_n709), .A3(new_n702), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n705), .B1(new_n710), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g510(.A(G50gat), .B1(new_n686), .B2(new_n341), .ZN(new_n712));
  INV_X1    g511(.A(new_n629), .ZN(new_n713));
  NOR4_X1   g512(.A1(new_n666), .A2(new_n713), .A3(G50gat), .A4(new_n341), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n572), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(KEYINPUT48), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n688), .A2(new_n342), .A3(new_n689), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n717), .A2(G50gat), .B1(new_n572), .B2(new_n714), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g518(.A1(new_n253), .A2(new_n608), .A3(new_n647), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT110), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n684), .A2(new_n571), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT111), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(KEYINPUT111), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n555), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g528(.A(new_n564), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(KEYINPUT112), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n735));
  INV_X1    g534(.A(G64gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n732), .A2(new_n735), .A3(new_n736), .A4(new_n733), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n741), .B2(new_n553), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n562), .A2(G71gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n742), .B(KEYINPUT50), .C1(new_n741), .C2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n726), .A2(new_n342), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g549(.A1(new_n253), .A2(new_n646), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT113), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n629), .A3(new_n722), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n609), .A2(G85gat), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n755), .A2(new_n727), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n676), .A2(new_n685), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n752), .A2(new_n608), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n578), .B1(new_n761), .B2(new_n727), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n757), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n757), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1336gat));
  NAND4_X1  g564(.A1(new_n755), .A2(new_n579), .A3(new_n490), .A4(new_n608), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n759), .A2(new_n760), .A3(new_n564), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n579), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT52), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n767), .A2(KEYINPUT115), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(KEYINPUT115), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(G92gat), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(new_n766), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(G1337gat));
  INV_X1    g574(.A(G99gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n608), .A2(new_n776), .A3(new_n561), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n755), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n759), .A2(new_n760), .A3(new_n553), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n776), .B2(new_n780), .ZN(G1338gat));
  NOR3_X1   g580(.A1(new_n609), .A2(G106gat), .A3(new_n341), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n755), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(G106gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n761), .B2(new_n342), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT53), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1339gat));
  INV_X1    g587(.A(new_n205), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n234), .A2(new_n236), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n243), .A2(new_n244), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT118), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n252), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n608), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n247), .A2(new_n252), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n596), .A2(new_n597), .A3(new_n574), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n605), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n603), .B1(new_n598), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n607), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n798), .B2(new_n800), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n796), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n678), .A2(new_n679), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n794), .A2(new_n804), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n678), .A2(new_n679), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n253), .A2(new_n609), .A3(new_n647), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n813), .A2(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(KEYINPUT117), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n812), .A2(new_n646), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n555), .A3(new_n569), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n564), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n351), .A2(new_n352), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n796), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n816), .A2(new_n342), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n564), .A2(new_n727), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n562), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n253), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n825), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n608), .A2(new_n344), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT119), .Z(new_n828));
  NAND2_X1  g627(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G120gat), .B1(new_n824), .B2(new_n609), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  NAND3_X1  g630(.A1(new_n818), .A2(new_n348), .A3(new_n645), .ZN(new_n832));
  OAI21_X1  g631(.A(G127gat), .B1(new_n824), .B2(new_n646), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n629), .A2(new_n564), .ZN(new_n835));
  AOI211_X1 g634(.A(G134gat), .B(new_n835), .C1(KEYINPUT120), .C2(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n817), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n629), .A3(new_n823), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(G134gat), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n841), .A2(new_n840), .A3(G134gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n810), .B1(new_n805), .B2(new_n795), .ZN(new_n845));
  AND4_X1   g644(.A1(new_n678), .A2(new_n794), .A3(new_n679), .A4(new_n804), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n646), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n814), .A2(new_n815), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n555), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n706), .A2(new_n341), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n253), .A2(G141gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n849), .A2(new_n564), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT122), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n706), .A2(new_n822), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n816), .B2(new_n341), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n806), .A2(new_n713), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n811), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n646), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n848), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n341), .A2(new_n858), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n265), .B1(new_n866), .B2(new_n796), .ZN(new_n867));
  INV_X1    g666(.A(new_n852), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n855), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n848), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n342), .ZN(new_n871));
  INV_X1    g670(.A(new_n864), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n862), .B2(new_n848), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n856), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n253), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n852), .A3(new_n854), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n869), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(new_n813), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n809), .A2(new_n629), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n880), .B2(new_n646), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n858), .B1(new_n881), .B2(new_n341), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n870), .A2(new_n864), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n856), .A2(new_n608), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT59), .B(G148gat), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n849), .A2(new_n564), .A3(new_n850), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT59), .B1(new_n887), .B2(new_n609), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n267), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n609), .A2(KEYINPUT59), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n886), .B(new_n889), .C1(new_n874), .C2(new_n890), .ZN(G1345gat));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n275), .B1(new_n866), .B2(new_n645), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n887), .A2(G155gat), .A3(new_n646), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G155gat), .B1(new_n874), .B2(new_n646), .ZN(new_n896));
  INV_X1    g695(.A(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(KEYINPUT123), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1346gat));
  NAND2_X1  g698(.A1(new_n849), .A2(new_n850), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(G162gat), .A3(new_n835), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT124), .ZN(new_n902));
  OAI21_X1  g701(.A(G162gat), .B1(new_n874), .B2(new_n807), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n564), .A2(new_n727), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n562), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n821), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n396), .A3(new_n253), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n816), .A2(new_n569), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n796), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(G1348gat));
  OAI21_X1  g711(.A(G176gat), .B1(new_n908), .B2(new_n609), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n397), .A3(new_n608), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  OAI21_X1  g714(.A(G183gat), .B1(new_n908), .B2(new_n646), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n910), .A2(new_n432), .A3(new_n645), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT60), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n429), .A3(new_n810), .ZN(new_n923));
  OAI21_X1  g722(.A(G190gat), .B1(new_n908), .B2(new_n713), .ZN(new_n924));
  XNOR2_X1  g723(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n924), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n706), .A2(new_n906), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n882), .B2(new_n883), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n796), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G197gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n253), .A2(G197gat), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n870), .A2(new_n850), .A3(new_n905), .A4(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT126), .Z(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n932), .B2(new_n796), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n937), .B(KEYINPUT126), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT127), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n939), .A2(new_n943), .ZN(G1352gat));
  NAND3_X1  g743(.A1(new_n870), .A2(new_n850), .A3(new_n905), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(G204gat), .A3(new_n609), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n608), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G204gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1353gat));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n645), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n953));
  INV_X1    g752(.A(G211gat), .ZN(new_n954));
  AOI211_X1 g753(.A(new_n953), .B(new_n954), .C1(new_n932), .C2(new_n645), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n645), .A2(new_n954), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n952), .A2(new_n955), .B1(new_n945), .B2(new_n956), .ZN(G1354gat));
  NAND2_X1  g756(.A1(new_n932), .A2(new_n629), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G218gat), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n807), .A2(G218gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n945), .B2(new_n960), .ZN(G1355gat));
endmodule


