//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G97), .A2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G77), .B2(G244), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G87), .A2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G58), .A2(G232), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n205), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AND2_X1   g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n203), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT1), .Z(new_n216));
  NOR2_X1   g0016(.A1(new_n203), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G20), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(new_n207), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(G1), .ZN(new_n243));
  OAI21_X1  g0043(.A(new_n243), .B1(G41), .B2(G45), .ZN(new_n244));
  INV_X1    g0044(.A(G274), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n244), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n208), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT66), .B(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G226), .ZN(new_n257));
  INV_X1    g0057(.A(G232), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n247), .B(new_n253), .C1(new_n262), .C2(new_n250), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n257), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n258), .A2(new_n259), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n254), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(new_n247), .A4(new_n253), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n264), .A2(G190), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n220), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT67), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n248), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT11), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n243), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT12), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n291), .B2(new_n207), .ZN(new_n295));
  INV_X1    g0095(.A(new_n278), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n289), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n293), .A2(new_n295), .B1(new_n207), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n276), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n264), .B2(new_n275), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n246), .B1(new_n271), .B2(new_n272), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n274), .B1(new_n304), .B2(new_n253), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n250), .B1(new_n270), .B2(new_n254), .ZN(new_n306));
  NOR4_X1   g0106(.A1(new_n306), .A2(KEYINPUT13), .A3(new_n246), .A4(new_n252), .ZN(new_n307));
  OAI21_X1  g0107(.A(G169), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n264), .A2(G179), .A3(new_n275), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n264), .A2(new_n275), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(G169), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n299), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n303), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n261), .B1(new_n208), .B2(new_n259), .C1(new_n256), .C2(new_n258), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n272), .C1(G107), .C2(new_n261), .ZN(new_n318));
  INV_X1    g0118(.A(new_n251), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G244), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n247), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT8), .B(G58), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT15), .B(G87), .Z(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n327), .B1(new_n329), .B2(new_n283), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n278), .B1(new_n284), .B2(new_n291), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n284), .B2(new_n297), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n316), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  INV_X1    g0135(.A(G222), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n261), .B1(new_n335), .B2(new_n259), .C1(new_n256), .C2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n272), .C1(G77), .C2(new_n261), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n247), .C1(new_n257), .C2(new_n251), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n339), .A2(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n280), .A2(G150), .ZN(new_n341));
  INV_X1    g0141(.A(G20), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n224), .A2(G50), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT8), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n223), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n223), .A2(KEYINPUT68), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G58), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n345), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n341), .B1(new_n342), .B2(new_n343), .C1(new_n350), .C2(new_n283), .ZN(new_n351));
  INV_X1    g0151(.A(G50), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n351), .A2(new_n279), .B1(new_n352), .B2(new_n291), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n296), .A2(KEYINPUT67), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT67), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n278), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n291), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(G50), .A3(new_n289), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n339), .A2(new_n323), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n340), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G190), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n339), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n353), .A2(KEYINPUT9), .A3(new_n358), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT10), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT9), .B1(new_n353), .B2(new_n358), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n339), .A2(G200), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n366), .A2(new_n367), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n370), .A3(new_n365), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT10), .B1(new_n372), .B2(new_n368), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n362), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G33), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT69), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT69), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n383), .A3(new_n342), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n261), .A2(G20), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(G68), .C1(new_n385), .C2(new_n379), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n346), .A2(new_n348), .A3(G68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n224), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n389), .A3(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n278), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n380), .A2(new_n382), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n342), .B2(new_n378), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT70), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n376), .B2(G33), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n248), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n377), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n379), .A2(G20), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(KEYINPUT71), .A3(new_n398), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n393), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n389), .B1(new_n403), .B2(new_n207), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n391), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n289), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT72), .B1(new_n350), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n346), .A2(new_n348), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT8), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n289), .A4(new_n345), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(new_n413), .A3(new_n357), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n350), .A2(new_n291), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n250), .A2(G232), .A3(new_n244), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n247), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n247), .A2(new_n418), .A3(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n265), .A2(new_n267), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n378), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n272), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n428), .A3(new_n363), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n256), .A2(new_n335), .B1(new_n257), .B2(new_n259), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n261), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n250), .B1(new_n431), .B2(new_n424), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n301), .B1(new_n432), .B2(new_n419), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n417), .A4(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n397), .A2(KEYINPUT71), .A3(new_n398), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT71), .B1(new_n397), .B2(new_n398), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(new_n385), .B2(new_n392), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G68), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT16), .B1(new_n439), .B2(new_n389), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n434), .B(new_n417), .C1(new_n440), .C2(new_n391), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n421), .A2(new_n422), .B1(new_n427), .B2(new_n272), .ZN(new_n445));
  INV_X1    g0245(.A(G179), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n430), .A2(new_n261), .B1(G33), .B2(G87), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n247), .B(new_n418), .C1(new_n447), .C2(new_n250), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n445), .A2(new_n446), .B1(new_n448), .B2(new_n323), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT18), .B(new_n449), .C1(new_n406), .C2(new_n416), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT74), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n406), .B2(new_n416), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n451), .A3(new_n454), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n444), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n321), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n332), .B1(G190), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n301), .B2(new_n459), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n334), .A2(new_n374), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n243), .A2(G33), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n357), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G107), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n291), .A2(new_n466), .ZN(new_n469));
  XOR2_X1   g0269(.A(new_n469), .B(KEYINPUT25), .Z(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT86), .A2(G87), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n375), .A2(new_n377), .A3(new_n471), .A4(new_n342), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT22), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n261), .A2(new_n474), .A3(new_n342), .A4(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n342), .A2(G33), .A3(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n466), .A2(G20), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT23), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n473), .B2(new_n475), .ZN(new_n484));
  INV_X1    g0284(.A(new_n482), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(new_n477), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n483), .A2(new_n486), .B1(KEYINPUT87), .B2(KEYINPUT24), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n468), .B(new_n470), .C1(new_n487), .C2(new_n296), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT77), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G41), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n249), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n245), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n243), .A2(G45), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT76), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n490), .A2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT76), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(new_n243), .A4(G45), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n493), .A2(new_n496), .A3(new_n250), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(G264), .A3(new_n250), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n375), .A2(new_n377), .A3(G257), .A4(G1698), .ZN(new_n505));
  OR2_X1    g0305(.A1(KEYINPUT88), .A2(G294), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT88), .A2(G294), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(G33), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n375), .A2(new_n377), .A3(G250), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n505), .B(new_n508), .C1(new_n509), .C2(new_n256), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n272), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n501), .A2(new_n504), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G169), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n504), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT89), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT89), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(new_n504), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n501), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n513), .B1(new_n518), .B2(new_n446), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n488), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n512), .A2(G190), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n518), .B2(new_n301), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n488), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n292), .A2(G97), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n465), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n466), .A2(KEYINPUT6), .A3(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n466), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n531), .B2(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n280), .A2(G77), .ZN(new_n534));
  XOR2_X1   g0334(.A(new_n534), .B(KEYINPUT75), .Z(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n535), .C1(new_n403), .C2(new_n466), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n527), .B1(new_n536), .B2(new_n278), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n425), .A2(new_n261), .A3(G244), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n425), .A2(new_n261), .A3(KEYINPUT4), .A4(G244), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n272), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n503), .A2(G257), .A3(new_n250), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(G190), .A3(new_n501), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT78), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n501), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n546), .B1(new_n544), .B2(new_n272), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(KEYINPUT78), .A3(G190), .A4(new_n501), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n537), .A2(new_n550), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n323), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n446), .A3(new_n501), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n438), .A2(G107), .B1(G20), .B2(new_n532), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n296), .B1(new_n558), .B2(new_n535), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n556), .B(new_n557), .C1(new_n559), .C2(new_n527), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT19), .B1(new_n282), .B2(G97), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n342), .B1(new_n254), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n530), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n261), .A2(new_n342), .A3(G68), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT80), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n261), .A2(KEYINPUT80), .A3(new_n342), .A4(G68), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n278), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n329), .A2(new_n291), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n328), .B(KEYINPUT81), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n357), .A3(new_n464), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G244), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n256), .B2(new_n208), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(new_n261), .ZN(new_n579));
  INV_X1    g0379(.A(G116), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n272), .B1(new_n248), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(G274), .B1(KEYINPUT79), .B2(G250), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n250), .B1(new_n495), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n495), .A2(new_n584), .A3(G250), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n579), .A2(new_n581), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n446), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n581), .B1(new_n578), .B2(new_n261), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n583), .A2(new_n586), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n323), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n576), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n465), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(G200), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n571), .A2(new_n278), .B1(new_n291), .B2(new_n329), .ZN(new_n597));
  OAI21_X1  g0397(.A(G190), .B1(new_n589), .B2(new_n590), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n555), .A2(new_n560), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n523), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n375), .A2(new_n377), .A3(G257), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n256), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n425), .A2(new_n261), .A3(KEYINPUT82), .A4(G257), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n378), .A2(G303), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n261), .A2(G264), .A3(G1698), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n272), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n503), .A2(G270), .A3(new_n250), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n501), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n543), .B(new_n342), .C1(G33), .C2(new_n526), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n580), .A2(G20), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT83), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n613), .A2(new_n278), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n615), .A2(KEYINPUT83), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n291), .A2(new_n278), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n580), .B1(new_n243), .B2(G33), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n620), .A2(new_n621), .B1(new_n580), .B2(new_n291), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n323), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n612), .A2(new_n623), .A3(KEYINPUT21), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT21), .B1(new_n612), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n622), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n500), .B1(new_n609), .B2(new_n272), .ZN(new_n628));
  AND4_X1   g0428(.A1(G179), .A2(new_n627), .A3(new_n611), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n612), .A2(G200), .ZN(new_n632));
  INV_X1    g0432(.A(new_n627), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(KEYINPUT84), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n301), .B1(new_n628), .B2(new_n611), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n627), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n628), .A2(G190), .A3(new_n611), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT85), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n637), .A3(new_n641), .A4(new_n638), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n463), .A2(new_n602), .A3(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n455), .A2(new_n450), .ZN(new_n645));
  INV_X1    g0445(.A(new_n303), .ZN(new_n646));
  INV_X1    g0446(.A(new_n333), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n646), .A2(new_n647), .B1(new_n314), .B2(new_n315), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(new_n444), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n371), .A2(new_n373), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n362), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n593), .A2(new_n599), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n560), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n536), .A2(new_n278), .ZN(new_n655));
  INV_X1    g0455(.A(new_n527), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n655), .A2(new_n656), .B1(new_n323), .B2(new_n551), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n600), .A2(new_n657), .A3(KEYINPUT26), .A4(new_n557), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n470), .ZN(new_n660));
  NAND2_X1  g0460(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n481), .A2(new_n482), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n485), .B1(new_n484), .B2(new_n477), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI211_X1 g0464(.A(new_n467), .B(new_n660), .C1(new_n664), .C2(new_n278), .ZN(new_n665));
  INV_X1    g0465(.A(new_n522), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n488), .A2(new_n519), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n631), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n659), .B(new_n593), .C1(new_n669), .C2(new_n601), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n651), .B1(new_n462), .B2(new_n671), .ZN(G369));
  NOR2_X1   g0472(.A1(new_n290), .A2(G20), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n243), .ZN(new_n674));
  XNOR2_X1  g0474(.A(KEYINPUT90), .B(KEYINPUT27), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n627), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT92), .Z(new_n683));
  NOR3_X1   g0483(.A1(new_n624), .A2(new_n629), .A3(new_n625), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n643), .B2(new_n683), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT93), .B(G330), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n681), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n667), .B(new_n520), .C1(new_n665), .C2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n668), .A2(new_n681), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n684), .A2(new_n520), .B1(new_n665), .B2(new_n666), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n690), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n217), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n565), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n225), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT94), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(new_n593), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n555), .A2(new_n560), .A3(new_n600), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n696), .B2(new_n708), .ZN(new_n709));
  AOI211_X1 g0509(.A(KEYINPUT29), .B(new_n681), .C1(new_n709), .C2(new_n659), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n670), .B2(new_n690), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n628), .A2(new_n587), .A3(G179), .A4(new_n611), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n511), .A2(new_n504), .A3(new_n516), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n516), .B1(new_n511), .B2(new_n504), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n716), .A2(new_n717), .A3(new_n500), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n715), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n553), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n553), .A2(new_n515), .A3(new_n501), .A4(new_n517), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n714), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n587), .B1(new_n628), .B2(new_n611), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n518), .A2(new_n723), .A3(new_n446), .A4(new_n551), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n681), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT95), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n681), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT95), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n602), .A2(new_n643), .A3(new_n690), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n728), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(new_n688), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n713), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n706), .B1(new_n738), .B2(G1), .ZN(G364));
  AOI21_X1  g0539(.A(new_n220), .B1(G20), .B2(new_n323), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n342), .A2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n301), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n741), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(G329), .B1(G283), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT99), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n342), .A2(new_n363), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n446), .A2(new_n301), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G326), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n755), .A2(new_n741), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  OAI22_X1  g0561(.A1(new_n757), .A2(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n754), .A2(new_n749), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n261), .B(new_n762), .C1(G303), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n753), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n446), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(G322), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n767), .A2(new_n741), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n506), .A2(new_n507), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n342), .B1(new_n742), .B2(G190), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n770), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT100), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n743), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT32), .Z(new_n779));
  OAI221_X1 g0579(.A(new_n261), .B1(new_n772), .B2(new_n284), .C1(new_n466), .C2(new_n750), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n764), .A2(G87), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n207), .B2(new_n760), .ZN(new_n782));
  INV_X1    g0582(.A(new_n774), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n780), .B(new_n782), .C1(G97), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n769), .A2(new_n410), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n779), .B(new_n786), .C1(G50), .C2(new_n756), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n740), .B1(new_n776), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n740), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n699), .A2(new_n261), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G45), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n238), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n225), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n796), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n261), .A2(G355), .A3(new_n217), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G116), .B2(new_n217), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT97), .Z(new_n801));
  OAI21_X1  g0601(.A(new_n792), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n673), .A2(G45), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT96), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT96), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(G1), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n700), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n686), .A2(new_n791), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n788), .A2(new_n802), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n687), .A2(new_n688), .ZN(new_n810));
  INV_X1    g0610(.A(new_n807), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n689), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(new_n812), .ZN(G396));
  NOR2_X1   g0613(.A1(new_n333), .A2(new_n681), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n681), .A2(new_n332), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n461), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n814), .B1(new_n816), .B2(new_n333), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(new_n790), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n740), .A2(new_n789), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n284), .ZN(new_n821));
  INV_X1    g0621(.A(new_n772), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G143), .A2(new_n769), .B1(new_n822), .B2(G159), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n757), .C1(new_n825), .C2(new_n760), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n748), .A2(G132), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G50), .A2(new_n764), .B1(new_n751), .B2(G68), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n827), .A2(new_n261), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n410), .B2(new_n783), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n748), .A2(G311), .B1(G97), .B2(new_n783), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n751), .A2(G87), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n760), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n763), .A2(new_n466), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n768), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G303), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n378), .B1(new_n580), .B2(new_n772), .C1(new_n757), .C2(new_n839), .ZN(new_n840));
  NOR4_X1   g0640(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n740), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n818), .A2(new_n807), .A3(new_n821), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n681), .B1(new_n709), .B2(new_n659), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(new_n817), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(new_n737), .Z(new_n846));
  OAI21_X1  g0646(.A(new_n843), .B1(new_n846), .B2(new_n807), .ZN(G384));
  AOI21_X1  g0647(.A(new_n312), .B1(new_n311), .B2(G169), .ZN(new_n848));
  AOI211_X1 g0648(.A(KEYINPUT14), .B(new_n323), .C1(new_n264), .C2(new_n275), .ZN(new_n849));
  INV_X1    g0649(.A(new_n310), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n315), .A2(new_n681), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n646), .B(new_n852), .C1(new_n851), .C2(new_n299), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n817), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n726), .A2(new_n727), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n735), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT106), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n679), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n406), .A2(new_n416), .B1(new_n449), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n441), .ZN(new_n865));
  INV_X1    g0665(.A(new_n441), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n386), .A2(new_n389), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n405), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n279), .A3(new_n390), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT104), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n869), .A2(new_n417), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n869), .B2(new_n417), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n449), .A2(new_n862), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n866), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n865), .B1(new_n875), .B2(new_n864), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n862), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n458), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT38), .B(new_n876), .C1(new_n458), .C2(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n316), .B2(new_n852), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n856), .B1(new_n884), .B2(new_n853), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n735), .A2(new_n859), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n817), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n861), .A2(new_n882), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n862), .B1(new_n406), .B2(new_n416), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n435), .A2(new_n443), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n645), .ZN(new_n893));
  INV_X1    g0693(.A(new_n865), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n864), .B1(new_n863), .B2(new_n441), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n879), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n881), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n885), .A2(new_n886), .A3(new_n817), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT40), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n890), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n463), .A2(new_n886), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n688), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n463), .B1(new_n710), .B2(new_n712), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n651), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT105), .Z(new_n908));
  XNOR2_X1  g0708(.A(new_n905), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n880), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n898), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n851), .A2(new_n299), .A3(new_n681), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n670), .A2(new_n690), .A3(new_n817), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n814), .B(KEYINPUT102), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n882), .A2(new_n885), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n455), .A2(new_n450), .A3(new_n679), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n909), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n243), .B2(new_n673), .ZN(new_n922));
  OAI211_X1 g0722(.A(G20), .B(new_n221), .C1(new_n532), .C2(KEYINPUT35), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n580), .B(new_n923), .C1(KEYINPUT35), .C2(new_n532), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  NAND3_X1  g0725(.A1(new_n797), .A2(G77), .A3(new_n387), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(G50), .B2(new_n207), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(G1), .A3(new_n290), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n922), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT107), .Z(G367));
  OAI211_X1 g0730(.A(new_n555), .B(new_n560), .C1(new_n537), .C2(new_n690), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT108), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n560), .B2(new_n690), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n694), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n595), .A2(new_n597), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n681), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n600), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n593), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT109), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n934), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n684), .A2(new_n681), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n933), .A2(new_n520), .A3(new_n667), .A4(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n560), .B1(new_n932), .B2(new_n520), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(new_n690), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n942), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n941), .B(new_n948), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n700), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n943), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n693), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT110), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n523), .B2(new_n952), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(KEYINPUT111), .A3(new_n689), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n689), .A2(KEYINPUT111), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n957), .B(new_n954), .C1(new_n523), .C2(new_n952), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n933), .A2(new_n697), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT45), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n932), .A2(new_n696), .A3(new_n690), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT44), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n694), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n695), .A3(new_n963), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n965), .A3(new_n738), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n951), .B1(new_n967), .B2(new_n738), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n949), .B1(new_n968), .B2(new_n806), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n750), .A2(new_n284), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G159), .B2(new_n759), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n349), .B2(new_n763), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n756), .A2(G143), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n772), .A2(new_n352), .B1(new_n743), .B2(new_n824), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n972), .A2(new_n378), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n207), .B2(new_n774), .C1(new_n825), .C2(new_n768), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n760), .A2(new_n773), .B1(new_n839), .B2(new_n768), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n763), .A2(new_n580), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(G311), .C2(new_n756), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n378), .B1(new_n743), .B2(new_n981), .C1(new_n526), .C2(new_n750), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT113), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n980), .B(new_n983), .C1(new_n834), .C2(new_n772), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n774), .A2(new_n466), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n740), .ZN(new_n988));
  INV_X1    g0788(.A(new_n791), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n938), .A2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n792), .B1(new_n217), .B2(new_n329), .C1(new_n230), .C2(new_n794), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT112), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n988), .A2(new_n807), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n969), .A2(new_n993), .ZN(G387));
  NAND2_X1  g0794(.A1(new_n956), .A2(new_n958), .ZN(new_n995));
  INV_X1    g0795(.A(new_n738), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n701), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n996), .B2(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n326), .A2(new_n352), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT50), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n207), .A2(new_n284), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n702), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n1000), .A2(G45), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n793), .B1(new_n234), .B2(new_n795), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n217), .A3(new_n261), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n217), .A2(G107), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n792), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n693), .A2(new_n791), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n768), .A2(new_n352), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n760), .A2(new_n350), .B1(new_n825), .B2(new_n743), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n574), .C2(new_n783), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n764), .A2(G77), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n757), .A2(new_n777), .B1(new_n750), .B2(new_n526), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G68), .B2(new_n822), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n261), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G322), .A2(new_n756), .B1(new_n759), .B2(G311), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n839), .B2(new_n772), .C1(new_n981), .C2(new_n768), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT48), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n834), .B2(new_n774), .C1(new_n773), .C2(new_n763), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT114), .Z(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT49), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n378), .B1(new_n743), .B2(new_n758), .C1(new_n580), .C2(new_n750), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT115), .Z(new_n1024));
  OAI21_X1  g0824(.A(new_n1016), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n811), .B(new_n1009), .C1(new_n1025), .C2(new_n740), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n959), .A2(new_n806), .B1(new_n1008), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n998), .A2(new_n1027), .ZN(G393));
  AND2_X1   g0828(.A1(new_n965), .A2(new_n966), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n738), .B2(new_n959), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n701), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n967), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n806), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n792), .B1(new_n526), .B2(new_n217), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n241), .B2(new_n793), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n769), .A2(G311), .B1(new_n756), .B2(G317), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n261), .B1(new_n744), .B2(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n466), .B2(new_n750), .C1(new_n834), .C2(new_n763), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT116), .Z(new_n1040));
  AOI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(G303), .C2(new_n759), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n580), .B2(new_n774), .C1(new_n837), .C2(new_n772), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT117), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n760), .A2(new_n352), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n769), .A2(G159), .B1(new_n756), .B2(G150), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n833), .B1(new_n207), .B2(new_n763), .C1(new_n325), .C2(new_n772), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n378), .B1(new_n744), .B2(G143), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n783), .A2(G77), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n811), .B(new_n1035), .C1(new_n1052), .C2(new_n740), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n989), .B2(new_n933), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1032), .A2(new_n1033), .A3(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n910), .A2(new_n912), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n789), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n820), .A2(new_n350), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n781), .B(new_n1050), .C1(new_n466), .C2(new_n760), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n757), .A2(new_n834), .B1(new_n750), .B2(new_n207), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n378), .B1(new_n772), .B2(new_n526), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n580), .B2(new_n768), .C1(new_n837), .C2(new_n747), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n764), .A2(G150), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT53), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n378), .B(new_n1065), .C1(G125), .C2(new_n748), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n759), .A2(G137), .B1(new_n783), .B2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT54), .B(G143), .Z(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n772), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT120), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(G128), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1072), .B1(new_n352), .B2(new_n750), .C1(new_n1073), .C2(new_n757), .ZN(new_n1074));
  INV_X1    g0874(.A(G132), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n768), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1063), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n740), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1057), .A2(new_n807), .A3(new_n1058), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n913), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n916), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n844), .B2(new_n817), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n885), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1056), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n885), .A2(KEYINPUT118), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT118), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1087), .B(new_n856), .C1(new_n884), .C2(new_n853), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n917), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n1080), .A3(new_n898), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n736), .A2(new_n688), .A3(new_n885), .A4(new_n817), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1085), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n885), .A2(new_n886), .A3(G330), .A4(new_n817), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1090), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n917), .A2(new_n885), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(new_n1080), .B1(new_n910), .B2(new_n912), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT119), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1085), .A2(new_n1090), .A3(new_n1100), .A4(new_n1091), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n806), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1079), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(G330), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n906), .B(new_n651), .C1(new_n1105), .C2(new_n903), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n736), .A2(new_n688), .A3(new_n817), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1083), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1094), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n917), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n886), .A2(G330), .A3(new_n817), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1082), .B(new_n1091), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1106), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1093), .A2(new_n1114), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1115), .A2(new_n700), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1106), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1102), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1104), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(G378));
  INV_X1    g0922(.A(KEYINPUT57), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1106), .B(KEYINPUT123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1115), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n650), .A2(new_n361), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1127), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n374), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n862), .A2(new_n359), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n359), .A3(new_n862), .A4(new_n1130), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n882), .A2(new_n889), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n898), .A2(new_n817), .A3(new_n885), .A4(new_n886), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1136), .A2(new_n861), .B1(KEYINPUT40), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1138), .B2(new_n1105), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n920), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1135), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n902), .A2(G330), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n902), .B2(G330), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1105), .B(new_n1135), .C1(new_n890), .C2(new_n901), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n920), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1123), .B1(new_n1125), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1146), .A3(KEYINPUT57), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT124), .B1(new_n1125), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT124), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1115), .A2(new_n1124), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT57), .A4(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1148), .A2(new_n1150), .A3(new_n700), .A4(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1013), .B(new_n249), .C1(new_n207), .C2(new_n774), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n261), .B1(new_n748), .B2(G283), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n466), .B2(new_n768), .C1(new_n580), .C2(new_n757), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(new_n410), .C2(new_n751), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n574), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1159), .B1(new_n526), .B2(new_n760), .C1(new_n1160), .C2(new_n772), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT58), .Z(new_n1162));
  AOI22_X1  g0962(.A1(G128), .A2(new_n769), .B1(new_n822), .B2(G137), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n764), .A2(new_n1068), .B1(new_n783), .B2(G150), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n756), .A2(G125), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G132), .B2(new_n759), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G41), .B1(new_n744), .B2(G124), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n248), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G159), .B2(new_n751), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1168), .B2(new_n1167), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(G50), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n740), .B1(new_n1162), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n811), .B1(new_n352), .B2(new_n819), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT121), .Z(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(new_n1135), .C2(new_n790), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT122), .Z(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1151), .B2(new_n806), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1181), .ZN(G375));
  NAND3_X1  g0982(.A1(new_n1110), .A2(new_n1106), .A3(new_n1113), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1119), .A2(new_n950), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1111), .A2(new_n790), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n740), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1160), .A2(new_n774), .B1(new_n837), .B2(new_n757), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n970), .B(new_n1187), .C1(G303), .C2(new_n748), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n759), .A2(G116), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n822), .A2(G107), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n526), .A2(new_n763), .B1(new_n768), .B2(new_n834), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n261), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n261), .B1(new_n747), .B2(new_n1073), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n774), .A2(new_n352), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n760), .A2(new_n1069), .B1(new_n349), .B2(new_n750), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n763), .A2(new_n777), .B1(new_n772), .B2(new_n825), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n1075), .B2(new_n757), .C1(new_n824), .C2(new_n768), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1186), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1185), .A2(new_n811), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n820), .A2(new_n207), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n806), .A2(new_n1117), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1184), .A2(new_n1203), .ZN(G381));
  XNOR2_X1  g1004(.A(G375), .B(KEYINPUT125), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G378), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(G390), .A2(G396), .A3(G387), .A4(G393), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(G381), .A2(G384), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(G407));
  INV_X1    g1009(.A(G213), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1206), .B2(new_n680), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(G407), .ZN(G409));
  INV_X1    g1012(.A(G390), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT126), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n969), .B2(new_n993), .ZN(new_n1215));
  INV_X1    g1015(.A(G396), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n998), .A2(new_n1216), .A3(new_n1027), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n998), .B2(new_n1027), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1217), .C1(new_n969), .C2(new_n993), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1213), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G387), .A2(new_n1219), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G390), .B(new_n1223), .C1(new_n1219), .C2(new_n1215), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1210), .A2(G343), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1119), .B(new_n700), .C1(new_n1227), .C2(new_n1183), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1183), .A2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1203), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(G384), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1155), .A2(G378), .A3(new_n1181), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n806), .B1(new_n1153), .B2(new_n950), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1179), .B1(new_n1234), .B2(new_n1147), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1121), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1226), .B(new_n1232), .C1(new_n1233), .C2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1226), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1226), .A2(G2897), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1231), .B(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1237), .A2(new_n1238), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1226), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1238), .A3(new_n1244), .A4(new_n1231), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1225), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1237), .A2(KEYINPUT63), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1241), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1249), .B(new_n1250), .C1(new_n1254), .C2(new_n1237), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1248), .A2(new_n1255), .ZN(G405));
  NAND2_X1  g1056(.A1(G375), .A2(new_n1121), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1233), .A2(new_n1259), .A3(new_n1231), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1231), .B1(new_n1233), .B2(new_n1259), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1233), .A2(new_n1259), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1232), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1233), .A2(new_n1259), .A3(new_n1231), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1257), .A3(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1262), .A2(new_n1266), .A3(new_n1225), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1225), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G402));
endmodule


