//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n209), .B(new_n222), .C1(new_n226), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G50), .B(G68), .Z(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G97), .B(G107), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G223), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(G1698), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n251), .B1(new_n252), .B2(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G274), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n257), .A2(new_n261), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n265), .B2(G226), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G200), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n223), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT65), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(KEYINPUT65), .A3(new_n223), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n216), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT8), .B1(new_n216), .B2(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n281), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n276), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n286), .A3(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n202), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n279), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n267), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G190), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n269), .A2(new_n270), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n294), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n302), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n270), .A2(new_n295), .A3(new_n297), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n269), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n293), .B1(new_n296), .B2(G169), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n267), .A2(G179), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n287), .A2(new_n252), .B1(new_n286), .B2(G68), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n314), .A2(new_n315), .B1(G50), .B2(new_n280), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n315), .B2(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n276), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT11), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(KEYINPUT11), .A3(new_n276), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n291), .A2(new_n218), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT12), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(KEYINPUT12), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n278), .A2(G68), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n250), .A2(KEYINPUT72), .A3(G226), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT72), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n253), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n332), .B1(new_n334), .B2(new_n211), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n249), .A2(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G232), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n331), .A2(new_n335), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n257), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n262), .B1(new_n264), .B2(new_n219), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n330), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AOI211_X1 g0143(.A(KEYINPUT13), .B(new_n341), .C1(new_n339), .C2(new_n257), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n328), .B1(new_n329), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NOR4_X1   g0147(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT73), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n345), .B2(G190), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n346), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n352));
  OAI211_X1 g0152(.A(G169), .B(new_n352), .C1(new_n343), .C2(new_n344), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n340), .A2(new_n342), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n340), .A2(new_n330), .A3(new_n342), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(G179), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT76), .B(KEYINPUT14), .Z(new_n360));
  OAI211_X1 g0160(.A(new_n353), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n362));
  INV_X1    g0162(.A(new_n360), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n345), .B2(new_n358), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n353), .A4(new_n357), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n328), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n337), .A2(G238), .B1(G107), .B2(new_n249), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n250), .A2(G232), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT67), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n257), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n263), .B1(new_n265), .B2(G244), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(KEYINPUT68), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT68), .B1(new_n374), .B2(new_n375), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n358), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n377), .B2(new_n378), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT8), .B(G58), .Z(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n287), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(new_n276), .B1(new_n252), .B2(new_n291), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n278), .A2(G77), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n380), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n378), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(G200), .A3(new_n376), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n389), .B(KEYINPUT69), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n379), .C2(new_n347), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n313), .A2(new_n351), .A3(new_n367), .A4(new_n395), .ZN(new_n396));
  MUX2_X1   g0196(.A(new_n291), .B(new_n278), .S(new_n284), .Z(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n216), .A2(new_n218), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n280), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n247), .A2(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT7), .B(new_n286), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT78), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n249), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n286), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n253), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n399), .B(new_n403), .C1(new_n412), .C2(G68), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n406), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n403), .B1(new_n414), .B2(G68), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n276), .B1(new_n415), .B2(KEYINPUT16), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n398), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n276), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT7), .B1(new_n249), .B2(new_n286), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n410), .B(G20), .C1(new_n246), .C2(new_n248), .ZN(new_n420));
  OAI21_X1  g0220(.A(G68), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n403), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n423), .B2(new_n399), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n412), .A2(G68), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT16), .A3(new_n422), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT79), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n397), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n262), .B1(new_n264), .B2(new_n217), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n431), .B1(new_n255), .B2(new_n211), .C1(new_n254), .C2(new_n334), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n432), .B2(new_n257), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(new_n329), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(G190), .B2(new_n433), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n429), .B1(new_n428), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n397), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n413), .A2(new_n416), .A3(new_n398), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT79), .B1(new_n424), .B2(new_n426), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n433), .A2(new_n358), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n381), .B(new_n430), .C1(new_n432), .C2(new_n257), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT18), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(KEYINPUT18), .A3(new_n446), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n417), .A2(new_n427), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n445), .B1(new_n451), .B2(new_n439), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(KEYINPUT80), .A3(KEYINPUT18), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n438), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n396), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT21), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n286), .C1(G33), .C2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n272), .C1(new_n286), .C2(G116), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  OR3_X1    g0262(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT84), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n462), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n291), .B1(new_n277), .B2(G33), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n418), .A2(G116), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n291), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n249), .A2(G303), .ZN(new_n472));
  INV_X1    g0272(.A(G264), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n255), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G257), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n334), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n257), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n277), .B(G45), .C1(new_n478), .C2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(G274), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n479), .A2(new_n481), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n257), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n484), .B2(G270), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G169), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n457), .B1(new_n471), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(KEYINPUT21), .A3(G169), .A4(new_n486), .ZN(new_n490));
  INV_X1    g0290(.A(new_n486), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(G179), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n418), .A2(new_n467), .ZN(new_n494));
  INV_X1    g0294(.A(G107), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n291), .A2(new_n495), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n495), .A2(KEYINPUT23), .A3(G20), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT23), .B1(new_n495), .B2(G20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n501), .A2(new_n502), .B1(G20), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n253), .A2(new_n286), .A3(G87), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT22), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(KEYINPUT22), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n253), .A2(new_n286), .A3(G87), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT86), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n507), .A2(new_n509), .ZN(new_n514));
  OAI211_X1 g0314(.A(KEYINPUT87), .B(KEYINPUT24), .C1(new_n514), .C2(new_n504), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT86), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(new_n516), .A3(new_n511), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT87), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(new_n515), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n500), .B1(new_n520), .B2(new_n276), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G294), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n255), .B2(new_n475), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n334), .A2(new_n213), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n257), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n482), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n484), .A2(G264), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(G179), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n358), .B2(new_n529), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n493), .B1(new_n522), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n529), .A2(new_n347), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(G200), .B2(new_n529), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n486), .A2(new_n347), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G200), .B2(new_n486), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n521), .A2(new_n534), .B1(new_n471), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n495), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  INV_X1    g0338(.A(new_n242), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(KEYINPUT6), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n414), .A2(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n418), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n291), .A2(new_n459), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n494), .B2(new_n459), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n253), .A2(G244), .A3(new_n333), .ZN(new_n548));
  NOR2_X1   g0348(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n458), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n257), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n482), .B1(new_n484), .B2(G257), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT82), .B1(new_n554), .B2(G179), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n556), .A3(new_n381), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n358), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n546), .A2(new_n555), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n253), .A2(G238), .A3(new_n333), .ZN(new_n560));
  INV_X1    g0360(.A(G244), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n503), .C1(new_n255), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n257), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n260), .A2(G1), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n257), .A2(new_n213), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(G274), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G169), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n381), .C2(new_n567), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n253), .A2(new_n286), .A3(G68), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n286), .B1(new_n336), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n212), .A2(new_n459), .A3(new_n495), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n287), .B2(new_n459), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n276), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n385), .A2(new_n291), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n494), .C2(new_n385), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n563), .A2(G179), .A3(new_n566), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n358), .B1(new_n563), .B2(new_n566), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT83), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n570), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n543), .A2(new_n545), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n554), .A2(G200), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n347), .C2(new_n554), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n567), .A2(G200), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n418), .A2(G87), .A3(new_n467), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n578), .A3(new_n579), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n588), .B(new_n591), .C1(new_n347), .C2(new_n567), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n559), .A2(new_n584), .A3(new_n587), .A4(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n456), .A2(new_n532), .A3(new_n537), .A4(new_n593), .ZN(G372));
  NAND2_X1  g0394(.A1(new_n532), .A2(KEYINPUT88), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n559), .A2(new_n587), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n521), .A2(new_n534), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT88), .ZN(new_n602));
  INV_X1    g0402(.A(new_n531), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n521), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n604), .B2(new_n493), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n595), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n557), .A2(new_n546), .A3(new_n555), .A4(new_n558), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n599), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n598), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n592), .A3(new_n584), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(KEYINPUT26), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n456), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n436), .A2(new_n437), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n351), .A2(new_n390), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(new_n367), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT18), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n428), .B2(new_n445), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n449), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n311), .B1(new_n621), .B2(new_n308), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n622), .ZN(G369));
  NAND2_X1  g0423(.A1(new_n522), .A2(new_n531), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n290), .A2(G20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n277), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n631), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n597), .B1(new_n521), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n632), .B1(new_n624), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n493), .A2(new_n633), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n471), .A2(new_n633), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n493), .A2(new_n639), .B1(new_n471), .B2(new_n536), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n493), .B2(new_n639), .ZN(new_n641));
  INV_X1    g0441(.A(G330), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(G399));
  INV_X1    g0447(.A(new_n207), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(G41), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n574), .A2(G116), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G1), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n227), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT28), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n532), .A2(new_n593), .A3(new_n537), .A4(new_n633), .ZN(new_n655));
  XNOR2_X1  g0455(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n486), .B2(new_n381), .ZN(new_n658));
  INV_X1    g0458(.A(new_n554), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT90), .A4(G179), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n526), .A2(new_n563), .A3(new_n528), .A4(new_n566), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n491), .A2(G179), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n529), .A3(new_n554), .A4(new_n567), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n631), .B(new_n656), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n655), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n666), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT91), .B1(new_n662), .B2(new_n663), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n662), .A2(KEYINPUT91), .A3(new_n663), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n633), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(KEYINPUT31), .ZN(new_n676));
  OAI21_X1  g0476(.A(G330), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(KEYINPUT92), .B(G330), .C1(new_n670), .C2(new_n676), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n607), .A2(new_n599), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT26), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n684), .B(new_n598), .C1(KEYINPUT26), .C2(new_n611), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n600), .A2(new_n532), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT29), .B(new_n633), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n631), .B1(new_n606), .B2(new_n612), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n654), .B1(new_n691), .B2(G1), .ZN(G364));
  XNOR2_X1  g0492(.A(new_n625), .B(KEYINPUT93), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G45), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n649), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(G13), .A2(G33), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G20), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n641), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n286), .A2(G190), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n329), .A2(G179), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(G179), .A2(G200), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(G283), .A2(new_n705), .B1(new_n708), .B2(G329), .ZN(new_n709));
  INV_X1    g0509(.A(G322), .ZN(new_n710));
  NAND2_X1  g0510(.A1(G20), .A2(G190), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n711), .A2(new_n381), .A3(G200), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n709), .B(new_n249), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n381), .A2(new_n329), .ZN(new_n715));
  INV_X1    g0515(.A(new_n711), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n702), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(KEYINPUT33), .B(G317), .ZN(new_n721));
  AOI22_X1  g0521(.A1(G326), .A2(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G311), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n702), .A2(G179), .A3(new_n329), .ZN(new_n724));
  INV_X1    g0524(.A(G303), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n711), .A2(new_n329), .A3(G179), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT96), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n722), .B1(new_n723), .B2(new_n724), .C1(new_n725), .C2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n286), .B1(new_n706), .B2(G190), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n714), .B(new_n730), .C1(G294), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT97), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n719), .A2(new_n218), .B1(new_n704), .B2(new_n495), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n253), .B1(new_n731), .B2(new_n459), .C1(new_n717), .C2(new_n202), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(G58), .C2(new_n712), .ZN(new_n739));
  INV_X1    g0539(.A(G159), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n707), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT32), .ZN(new_n742));
  INV_X1    g0542(.A(new_n729), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G87), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G77), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n739), .A2(new_n742), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n735), .A2(new_n736), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n223), .B1(G20), .B2(new_n358), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n700), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n249), .A2(new_n207), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n228), .A2(new_n260), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n260), .C2(new_n240), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n648), .A2(new_n249), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(G355), .B1(new_n469), .B2(new_n648), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n697), .B1(new_n701), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n641), .B(new_n642), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n697), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT98), .ZN(G396));
  NOR2_X1   g0564(.A1(new_n390), .A2(new_n631), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n389), .A2(new_n631), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n394), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n390), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n682), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n679), .B2(new_n680), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n688), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n696), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(new_n688), .A3(new_n772), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n751), .A2(new_n698), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n697), .B1(new_n252), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n751), .ZN(new_n779));
  INV_X1    g0579(.A(new_n747), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n780), .A2(new_n469), .B1(new_n729), .B2(new_n495), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n705), .A2(G87), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n723), .B2(new_n707), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n713), .A2(new_n784), .B1(new_n719), .B2(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n249), .B1(new_n731), .B2(new_n459), .C1(new_n717), .C2(new_n725), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n781), .A2(new_n783), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n729), .A2(new_n202), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n704), .A2(new_n218), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n249), .B(new_n790), .C1(G132), .C2(new_n708), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n216), .B2(new_n731), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n718), .A2(G137), .B1(G143), .B2(new_n712), .ZN(new_n793));
  INV_X1    g0593(.A(G150), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n794), .B2(new_n719), .C1(new_n780), .C2(new_n740), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT34), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n789), .B(new_n792), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n788), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n778), .B1(new_n779), .B2(new_n799), .C1(new_n768), .C2(new_n699), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n776), .A2(new_n800), .ZN(G384));
  NAND2_X1  g0601(.A1(new_n362), .A2(new_n366), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n326), .B(KEYINPUT75), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n631), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n403), .B1(new_n412), .B2(G68), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n276), .B1(new_n807), .B2(KEYINPUT16), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT102), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(KEYINPUT102), .B(new_n276), .C1(new_n807), .C2(KEYINPUT16), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n426), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n629), .B1(new_n812), .B2(new_n439), .ZN(new_n813));
  AOI21_X1  g0613(.A(KEYINPUT80), .B1(new_n452), .B2(KEYINPUT18), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n428), .A2(new_n448), .A3(new_n618), .A4(new_n445), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n814), .A2(new_n815), .A3(new_n447), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n813), .B1(new_n816), .B2(new_n438), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT103), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n428), .A2(new_n435), .ZN(new_n819));
  INV_X1    g0619(.A(new_n629), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n443), .A2(new_n444), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n812), .B2(new_n439), .ZN(new_n822));
  OAI211_X1 g0622(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n819), .C2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT37), .B1(new_n819), .B2(new_n822), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT104), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n428), .A2(new_n821), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT37), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n824), .A2(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n817), .A2(new_n818), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(KEYINPUT103), .B(new_n813), .C1(new_n816), .C2(new_n438), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT38), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n824), .A2(new_n825), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n827), .A2(new_n828), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n823), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n813), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n449), .A2(new_n448), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(new_n453), .A3(new_n619), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n838), .B2(new_n615), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n839), .B2(KEYINPUT103), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n818), .B(new_n836), .C1(new_n838), .C2(new_n615), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT39), .B1(new_n832), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n818), .B1(new_n454), .B2(new_n836), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n831), .A4(new_n835), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT39), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n428), .B(new_n629), .C1(new_n615), .C2(new_n620), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n827), .B(KEYINPUT37), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n806), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(new_n846), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n767), .A2(new_n390), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n613), .A2(new_n633), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n765), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR3_X1    g0658(.A1(new_n328), .A2(KEYINPUT101), .A3(new_n633), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT101), .B1(new_n328), .B2(new_n633), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n351), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n804), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n328), .B(new_n633), .C1(new_n362), .C2(new_n366), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n854), .A2(new_n868), .B1(new_n620), .B2(new_n820), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n852), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n622), .B1(new_n455), .B2(new_n689), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n846), .A2(new_n850), .ZN(new_n874));
  INV_X1    g0674(.A(new_n656), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n672), .A2(new_n664), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n674), .A3(new_n666), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(new_n631), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT31), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(new_n655), .B1(new_n879), .B2(new_n675), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n367), .A2(new_n861), .A3(new_n351), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n880), .B(new_n768), .C1(new_n881), .C2(new_n865), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n873), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n867), .A2(new_n873), .A3(new_n768), .A4(new_n880), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n846), .B2(new_n853), .ZN(new_n886));
  OAI21_X1  g0686(.A(G330), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n880), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n642), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n455), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n882), .B1(new_n846), .B2(new_n850), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n854), .A2(new_n885), .B1(new_n893), .B2(new_n873), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n455), .A2(new_n888), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n887), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n872), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n872), .A2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n277), .B2(new_n693), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n900), .B2(new_n899), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n540), .B(KEYINPUT99), .Z(new_n903));
  INV_X1    g0703(.A(KEYINPUT35), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(G116), .A3(new_n226), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n906), .A2(KEYINPUT100), .B1(new_n904), .B2(new_n903), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(KEYINPUT100), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT36), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(KEYINPUT36), .ZN(new_n910));
  OAI21_X1  g0710(.A(G77), .B1(new_n216), .B2(new_n218), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n911), .A2(new_n227), .B1(G50), .B2(new_n218), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(G1), .A3(new_n290), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n902), .A2(new_n909), .A3(new_n910), .A4(new_n913), .ZN(G367));
  INV_X1    g0714(.A(KEYINPUT45), .ZN(new_n915));
  INV_X1    g0715(.A(new_n646), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n596), .B1(new_n585), .B2(new_n633), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n607), .A2(new_n631), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n915), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n646), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(KEYINPUT44), .A3(new_n920), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT44), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n646), .B2(new_n919), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n923), .A2(new_n927), .A3(new_n645), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n635), .A2(new_n636), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n637), .A2(new_n643), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n645), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n691), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n649), .B(KEYINPUT41), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n695), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n590), .A2(new_n631), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n599), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT106), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n599), .A2(KEYINPUT106), .A3(new_n935), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n938), .B(new_n939), .C1(new_n598), .C2(new_n935), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT107), .Z(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n604), .A2(new_n587), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n631), .B1(new_n944), .B2(new_n559), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n635), .A2(new_n596), .A3(new_n636), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n946), .B2(KEYINPUT42), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(new_n942), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n948), .A2(new_n947), .A3(new_n942), .A4(new_n941), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n644), .A2(new_n919), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(new_n952), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n941), .A2(new_n700), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n249), .B1(new_n719), .B2(new_n784), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT108), .B(G317), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G97), .A2(new_n705), .B1(new_n708), .B2(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n725), .B2(new_n713), .C1(new_n723), .C2(new_n717), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(G107), .C2(new_n732), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n785), .B2(new_n780), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n729), .A2(new_n469), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n704), .A2(new_n252), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n249), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT109), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n747), .A2(G50), .B1(new_n743), .B2(G58), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n732), .A2(G68), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G159), .A2(new_n720), .B1(new_n708), .B2(G137), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n718), .A2(G143), .B1(G150), .B2(new_n712), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n965), .A2(new_n967), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT47), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n779), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n977), .B2(new_n976), .ZN(new_n979));
  INV_X1    g0779(.A(new_n754), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n752), .B1(new_n207), .B2(new_n385), .C1(new_n980), .C2(new_n236), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n696), .A3(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n934), .A2(new_n958), .B1(new_n959), .B2(new_n982), .ZN(G387));
  AOI21_X1  g0783(.A(new_n253), .B1(new_n708), .B2(G326), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n469), .B2(new_n704), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n720), .A2(G311), .B1(new_n712), .B2(new_n961), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n710), .B2(new_n717), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G303), .B2(new_n747), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT48), .Z(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n785), .B2(new_n731), .C1(new_n784), .C2(new_n729), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT49), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n743), .A2(G77), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n794), .B2(new_n707), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n731), .A2(new_n385), .ZN(new_n997));
  INV_X1    g0797(.A(new_n724), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n998), .A2(G68), .B1(new_n712), .B2(G50), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n253), .C1(new_n459), .C2(new_n704), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n997), .B(new_n1000), .C1(new_n284), .C2(new_n720), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n717), .A2(new_n740), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT111), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n996), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n779), .B1(new_n993), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n980), .B1(new_n233), .B2(G45), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n651), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n757), .ZN(new_n1009));
  AOI21_X1  g0809(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n383), .A2(new_n202), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n651), .B(new_n1010), .C1(new_n1011), .C2(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(G107), .B2(new_n207), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n697), .B(new_n1006), .C1(new_n752), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT112), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OR3_X1    g0817(.A1(new_n635), .A2(G20), .A3(new_n699), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n931), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1017), .A2(new_n1018), .B1(new_n695), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n691), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n649), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n691), .A2(new_n1019), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G393));
  AOI21_X1  g0824(.A(new_n645), .B1(new_n923), .B2(new_n927), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n928), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n690), .A2(new_n931), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n923), .A2(new_n927), .A3(new_n645), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n650), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n923), .A2(new_n927), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n644), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n695), .A3(new_n1028), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n920), .A2(new_n700), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n747), .A2(new_n383), .B1(new_n743), .B2(G68), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n713), .A2(new_n740), .B1(new_n717), .B2(new_n794), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G50), .A2(new_n720), .B1(new_n708), .B2(G143), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n731), .A2(new_n252), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1040), .A2(new_n253), .A3(new_n782), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n718), .A2(G317), .B1(G311), .B2(new_n712), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n719), .A2(new_n725), .B1(new_n707), .B2(new_n710), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G294), .B2(new_n998), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n249), .B1(new_n704), .B2(new_n495), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G116), .B2(new_n732), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(new_n785), .C2(new_n729), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1039), .A2(new_n1043), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n751), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n752), .B1(new_n459), .B2(new_n207), .C1(new_n980), .C2(new_n243), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1034), .A2(new_n696), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1030), .A2(new_n1033), .A3(new_n1054), .ZN(G390));
  INV_X1    g0855(.A(KEYINPUT115), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n881), .A2(new_n865), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n769), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n889), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n771), .B2(new_n867), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1057), .B1(new_n890), .B2(new_n769), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n855), .B(new_n633), .C1(new_n685), .C2(new_n686), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n857), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n681), .B2(new_n1058), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1060), .A2(new_n858), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n871), .A2(new_n891), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n868), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n844), .B(new_n851), .C1(new_n805), .C2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n805), .B1(new_n1063), .B2(new_n867), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n874), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT114), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n874), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n681), .A2(new_n1058), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1059), .B1(new_n1079), .B2(new_n1070), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1056), .B(new_n1068), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1067), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1056), .B1(new_n1065), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1059), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n851), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n847), .B1(new_n853), .B2(new_n846), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n805), .B1(new_n858), .B2(new_n867), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1083), .A2(new_n1077), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1081), .A2(new_n649), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n697), .B1(new_n285), .B2(new_n777), .ZN(new_n1093));
  INV_X1    g0893(.A(G132), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n253), .B1(new_n731), .B2(new_n740), .C1(new_n713), .C2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G128), .A2(new_n718), .B1(new_n720), .B2(G137), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G50), .A2(new_n705), .B1(new_n708), .B2(G125), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  AOI211_X1 g0899(.A(new_n1095), .B(new_n1098), .C1(new_n747), .C2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n729), .A2(new_n794), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n720), .A2(G107), .B1(G116), .B2(new_n712), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n785), .B2(new_n717), .C1(new_n784), .C2(new_n707), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1104), .A2(new_n253), .A3(new_n790), .A4(new_n1041), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n747), .A2(G97), .B1(new_n743), .B2(G87), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1100), .A2(new_n1102), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1093), .B1(new_n1107), .B2(new_n779), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n698), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n695), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1092), .A2(new_n1112), .ZN(G378));
  INV_X1    g0913(.A(KEYINPUT118), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT55), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n313), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n293), .A2(new_n820), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n308), .A2(KEYINPUT55), .A3(new_n312), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1117), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT55), .B1(new_n308), .B2(new_n312), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1115), .B(new_n311), .C1(new_n303), .C2(new_n307), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1119), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1129), .B(G330), .C1(new_n884), .C2(new_n886), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n894), .B2(G330), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1114), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n870), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1129), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n887), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1130), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n620), .A2(new_n820), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n854), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n1069), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n805), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1114), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1090), .A2(new_n1077), .A3(new_n1066), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1067), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT57), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1142), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1136), .A2(new_n870), .A3(new_n1130), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(new_n1150), .A3(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n649), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1135), .A2(new_n698), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n718), .A2(G125), .B1(G128), .B2(new_n712), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n794), .B2(new_n731), .ZN(new_n1156));
  INV_X1    g0956(.A(G137), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n724), .A2(new_n1157), .B1(new_n719), .B2(new_n1094), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT116), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1156), .B(new_n1159), .C1(new_n743), .C2(new_n1099), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT59), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n245), .B(new_n259), .C1(new_n704), .C2(new_n740), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G124), .B2(new_n708), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n253), .A2(G41), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G50), .B(new_n1167), .C1(new_n245), .C2(new_n259), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n705), .A2(G58), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n712), .A2(G107), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n724), .A2(new_n385), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n994), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G97), .A2(new_n720), .B1(new_n708), .B2(G283), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n718), .A2(G116), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n972), .A3(new_n1167), .A4(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1168), .B1(new_n1176), .B2(KEYINPUT58), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1166), .B(new_n1177), .C1(KEYINPUT58), .C2(new_n1176), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n751), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n777), .A2(new_n202), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1154), .A2(new_n696), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1144), .B2(new_n695), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1153), .A2(new_n1183), .ZN(G375));
  NAND2_X1  g0984(.A1(new_n1065), .A2(new_n1082), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1068), .A2(new_n933), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n697), .B1(new_n218), .B2(new_n777), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n718), .A2(G294), .B1(G283), .B2(new_n712), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n469), .B2(new_n719), .C1(new_n725), .C2(new_n707), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1189), .A2(new_n253), .A3(new_n968), .A4(new_n997), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n747), .A2(G107), .B1(new_n743), .B2(G97), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n713), .A2(new_n1157), .B1(new_n717), .B2(new_n1094), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1169), .A2(new_n253), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G50), .C2(new_n732), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n720), .A2(new_n1099), .B1(new_n708), .B2(G128), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n794), .B2(new_n724), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G159), .B2(new_n743), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1190), .A2(new_n1191), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1187), .B1(new_n1198), .B2(new_n779), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1057), .B2(new_n698), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1066), .B2(new_n695), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1186), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT119), .ZN(G381));
  INV_X1    g1003(.A(G378), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1153), .A2(new_n1204), .A3(new_n1183), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1033), .A2(new_n1054), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n776), .A3(new_n800), .ZN(new_n1208));
  OR4_X1    g1008(.A1(G396), .A2(new_n1208), .A3(G387), .A4(G393), .ZN(new_n1209));
  OR3_X1    g1009(.A1(new_n1205), .A2(G381), .A3(new_n1209), .ZN(G407));
  OAI211_X1 g1010(.A(G407), .B(G213), .C1(G343), .C2(new_n1205), .ZN(G409));
  XNOR2_X1  g1011(.A(G393), .B(G396), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n959), .A2(new_n982), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n957), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n956), .B1(new_n951), .B2(new_n952), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n690), .B1(new_n1028), .B2(new_n1019), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n933), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G1), .B(new_n694), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1213), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT125), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1220), .A2(new_n1207), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G390), .B1(G387), .B2(KEYINPUT125), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1212), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT126), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT126), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1212), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT124), .B1(new_n1220), .B2(G390), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1220), .B2(G390), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1220), .A2(G390), .A3(KEYINPUT124), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  AOI221_X4 g1034(.A(KEYINPUT118), .B1(new_n1140), .B2(new_n1141), .C1(new_n1136), .C2(new_n1130), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1142), .B1(new_n1137), .B2(new_n1114), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1146), .B(new_n933), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT120), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT120), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1144), .A2(new_n1239), .A3(new_n933), .A4(new_n1146), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1136), .A2(new_n870), .A3(new_n1130), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1136), .A2(new_n1130), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n695), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1181), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1238), .A2(new_n1240), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1204), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1183), .C1(new_n1147), .C2(new_n1152), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT121), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n630), .A2(G213), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1252), .A3(new_n1248), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1185), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1065), .A2(new_n1082), .A3(KEYINPUT60), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1255), .A2(new_n1068), .A3(new_n649), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1201), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(G384), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .A4(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n630), .A2(G213), .A3(G2897), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1259), .B(new_n1263), .Z(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1248), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1244), .B1(KEYINPUT120), .B2(new_n1237), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1267), .B2(new_n1240), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1251), .B(new_n1259), .C1(new_n1266), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1228), .B(new_n1234), .C1(new_n1261), .C2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1274), .B2(new_n1260), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1253), .A2(new_n1251), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1252), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT122), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT122), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1250), .A2(new_n1280), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1281), .A3(new_n1264), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1276), .A2(new_n1282), .A3(KEYINPUT127), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT127), .B1(new_n1276), .B2(new_n1282), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1272), .B1(new_n1283), .B2(new_n1284), .ZN(G405));
  NAND2_X1  g1085(.A1(G375), .A2(G378), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1205), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1259), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1288), .B(new_n1289), .ZN(G402));
endmodule


