//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1220, new_n1221,
    new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT66), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n461), .A2(new_n464), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n470), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n476), .A2(G126), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  NAND2_X1  g069(.A1(G75), .A2(G543), .ZN(new_n495));
  XOR2_X1   g070(.A(KEYINPUT5), .B(G543), .Z(new_n496));
  INV_X1    g071(.A(G62), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(G50), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G166));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .A3(new_n512), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n517), .A3(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n507), .A2(new_n503), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n510), .A2(new_n520), .A3(new_n522), .A4(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n518), .A2(new_n528), .B1(new_n529), .B2(new_n523), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT72), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n509), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(new_n535), .B2(G651), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  AOI211_X1 g112(.A(KEYINPUT71), .B(new_n537), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n531), .B1(new_n536), .B2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n507), .B(KEYINPUT69), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n518), .A2(new_n547), .B1(new_n548), .B2(new_n523), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n545), .B(new_n546), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n549), .B(new_n550), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n546), .B1(new_n555), .B2(new_n545), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n496), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n524), .B2(G91), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n515), .A2(new_n517), .A3(G53), .A4(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n503), .B2(new_n511), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n570), .A2(new_n571), .A3(G53), .A4(new_n517), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n568), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n505), .B(new_n577), .ZN(G303));
  OAI21_X1  g153(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n519), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n524), .A2(G87), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n503), .A2(G48), .A3(G543), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n523), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n507), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n537), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n542), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n537), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n519), .A2(G47), .B1(new_n524), .B2(G85), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n599), .A2(KEYINPUT79), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT79), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  OR2_X1    g181(.A1(KEYINPUT80), .A2(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(KEYINPUT80), .A2(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(KEYINPUT81), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n613), .A2(new_n524), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n611), .C1(new_n523), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n519), .A2(G54), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n496), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n606), .B1(G868), .B2(new_n623), .ZN(G284));
  OAI21_X1  g199(.A(new_n606), .B1(G868), .B2(new_n623), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(new_n566), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n568), .A2(new_n572), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT75), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n626), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n623), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n623), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n557), .B2(G868), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n482), .A2(G135), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n477), .A2(G123), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n464), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n462), .A2(new_n468), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1341), .B(G1348), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2443), .B(G2446), .Z(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(G14), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n667), .ZN(G401));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(new_n678), .C1(new_n674), .C2(new_n676), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n674), .A3(new_n676), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT18), .Z(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n689), .A2(new_n694), .A3(new_n692), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n697));
  AOI211_X1 g272(.A(new_n693), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT89), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(G288), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT88), .B(G16), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1971), .Z(new_n717));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n592), .B2(G16), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n712), .B(new_n717), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n604), .A2(new_n714), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G24), .B2(new_n714), .ZN(new_n726));
  INV_X1    g301(.A(G1986), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n723), .A2(KEYINPUT34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n482), .A2(G131), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n464), .A2(G107), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n476), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G119), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n730), .B1(new_n731), .B2(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G25), .B(new_n736), .S(G29), .Z(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n729), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n728), .A2(KEYINPUT90), .A3(new_n740), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n724), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n724), .B(new_n748), .C1(new_n743), .C2(new_n744), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G140), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n464), .A2(G116), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G128), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n751), .B1(new_n752), .B2(new_n753), .C1(new_n734), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT92), .ZN(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n709), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n709), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n764), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n623), .B2(G16), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(G1348), .ZN(new_n771));
  INV_X1    g346(.A(new_n649), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n482), .A2(G139), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n464), .B2(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G33), .B(new_n782), .S(G29), .Z(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n770), .A2(G1348), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n768), .A2(new_n773), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n758), .A2(G35), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G162), .B2(new_n758), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT29), .Z(new_n789));
  INV_X1    g364(.A(G2090), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n474), .A2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT24), .ZN(new_n794));
  INV_X1    g369(.A(G34), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n792), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n793), .B1(new_n792), .B2(new_n797), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(G28), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n758), .B1(new_n800), .B2(G28), .ZN(new_n802));
  AND2_X1   g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n709), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n709), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n791), .A2(new_n798), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n482), .A2(G141), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n477), .A2(G129), .ZN(new_n814));
  NAND3_X1  g389(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT26), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n817), .A2(new_n818), .B1(G105), .B2(new_n468), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n813), .A2(new_n814), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n758), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n758), .B2(G32), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT27), .B(G1996), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n823), .A2(new_n824), .B1(new_n783), .B2(G2072), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n758), .A2(G27), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G164), .B2(new_n758), .ZN(new_n827));
  INV_X1    g402(.A(G2078), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n825), .B(new_n829), .C1(new_n823), .C2(new_n824), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n767), .A2(new_n786), .A3(new_n811), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n714), .A2(G19), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n557), .B2(new_n714), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G1341), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n713), .A2(G20), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT96), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT23), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n631), .B2(new_n709), .ZN(new_n838));
  INV_X1    g413(.A(G1956), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n789), .B2(new_n790), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n831), .B(new_n834), .C1(KEYINPUT97), .C2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n841), .A2(KEYINPUT97), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n750), .A2(new_n844), .ZN(G311));
  NAND2_X1  g420(.A1(new_n750), .A2(new_n844), .ZN(G150));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n518), .A2(new_n847), .B1(new_n848), .B2(new_n523), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n542), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n537), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  INV_X1    g434(.A(new_n856), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n554), .B2(new_n556), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n545), .A3(new_n555), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n623), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT99), .Z(new_n869));
  OAI21_X1  g444(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n859), .B1(new_n869), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n649), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n484), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n755), .B(new_n493), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(new_n782), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n820), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n482), .A2(G142), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n464), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n477), .B2(G130), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(new_n653), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n736), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n875), .B(new_n782), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n821), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n877), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n877), .A2(new_n886), .ZN(new_n890));
  INV_X1    g465(.A(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n889), .A2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n874), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n873), .A3(new_n887), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n631), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(G299), .A2(KEYINPUT101), .A3(new_n623), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n631), .A2(new_n902), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  AND3_X1   g485(.A1(G299), .A2(KEYINPUT101), .A3(new_n623), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT101), .B1(G299), .B2(new_n623), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n904), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n908), .B1(new_n915), .B2(KEYINPUT104), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  AOI211_X1 g492(.A(new_n917), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n863), .B(new_n636), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n904), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT102), .B1(new_n903), .B2(new_n904), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n906), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(KEYINPUT103), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n924), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G288), .B(new_n505), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n592), .B1(new_n602), .B2(new_n603), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n602), .A2(new_n592), .A3(new_n603), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n933), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n930), .A2(new_n931), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n921), .A2(new_n943), .A3(new_n925), .A4(new_n928), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n932), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n932), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g523(.A(new_n947), .B1(G868), .B2(new_n856), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  INV_X1    g526(.A(new_n909), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n924), .A2(new_n951), .B1(new_n905), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G301), .A2(G168), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n531), .B(G286), .C1(new_n536), .C2(new_n538), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n555), .A2(new_n545), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT74), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n856), .B1(new_n958), .B2(new_n553), .ZN(new_n959));
  INV_X1    g534(.A(new_n862), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n861), .A2(new_n862), .A3(new_n954), .A4(new_n955), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT107), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n906), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n913), .B2(new_n914), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n962), .B2(new_n961), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n952), .A2(new_n905), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n966), .B2(KEYINPUT41), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n961), .A2(new_n962), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n964), .A2(new_n968), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n941), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n952), .B1(new_n922), .B2(new_n923), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n917), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n908), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n967), .B1(new_n980), .B2(new_n971), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n941), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n950), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n907), .B1(new_n977), .B2(new_n917), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n963), .B1(new_n984), .B2(new_n979), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n975), .B1(new_n985), .B2(new_n967), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n971), .B1(new_n916), .B2(new_n918), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(new_n941), .A3(new_n968), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n989));
  AND4_X1   g564(.A1(new_n897), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT44), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n970), .A2(new_n971), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n967), .B1(new_n992), .B2(KEYINPUT107), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n941), .B1(new_n993), .B2(new_n973), .ZN(new_n994));
  INV_X1    g569(.A(new_n989), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G37), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n988), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT108), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n996), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n981), .B2(new_n941), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n976), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n988), .A2(new_n897), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n941), .B1(new_n987), .B2(new_n968), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n995), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n998), .A2(new_n1002), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n991), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n991), .B2(new_n1007), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n493), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT110), .B(G40), .Z(new_n1016));
  OR3_X1    g591(.A1(new_n465), .A2(new_n472), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n493), .A2(new_n1023), .A3(new_n1012), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1022), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(G1956), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n628), .A2(new_n566), .A3(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1030), .B(new_n1021), .C1(new_n1025), .C2(G1956), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1022), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1036), .A2(new_n1020), .B1(new_n1037), .B2(new_n839), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1348), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1022), .A2(new_n1018), .A3(KEYINPUT116), .A4(new_n1024), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1017), .A2(new_n1013), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n762), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT60), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n902), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(KEYINPUT60), .A3(new_n1048), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1040), .A2(new_n1041), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  INV_X1    g628(.A(G1996), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1015), .A2(new_n1018), .A3(new_n1054), .A4(new_n1019), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  AOI22_X1  g632(.A1(new_n1055), .A2(KEYINPUT117), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1036), .A2(new_n1059), .A3(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n557), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1053), .B1(new_n1062), .B2(KEYINPUT59), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n1064));
  INV_X1    g639(.A(new_n557), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(KEYINPUT119), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1063), .A2(new_n1064), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1032), .A2(new_n1072), .A3(KEYINPUT61), .A4(new_n1033), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1046), .A2(KEYINPUT60), .A3(new_n902), .A4(new_n1048), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1077), .B2(new_n1033), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1052), .A2(new_n1071), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n902), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1032), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1081), .A2(new_n1082), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT122), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1047), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT111), .B1(G288), .B2(new_n1090), .ZN(new_n1091));
  OR3_X1    g666(.A1(G288), .A2(KEYINPUT111), .A3(new_n1090), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1090), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1981), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n592), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT112), .B(G86), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n583), .B1(new_n523), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(G1981), .B1(new_n1100), .B2(new_n588), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT49), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(KEYINPUT49), .A3(new_n1101), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1089), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1094), .A2(new_n1096), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G303), .A2(G8), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1036), .A2(G1971), .B1(new_n1037), .B2(G2090), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(G8), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1111), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1108), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT125), .B(G1961), .Z(new_n1118));
  NAND3_X1  g693(.A1(new_n1043), .A2(new_n1045), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(G2078), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n828), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1123), .B(new_n465), .C1(new_n1124), .C2(new_n472), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n473), .A2(KEYINPUT126), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1015), .A2(new_n1125), .A3(new_n1019), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1036), .A2(KEYINPUT53), .A3(new_n828), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(new_n1130), .A3(new_n1122), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1129), .B(KEYINPUT54), .C1(G171), .C2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1128), .A2(G171), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(G171), .B2(new_n1131), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1117), .B(new_n1132), .C1(new_n1134), .C2(KEYINPUT54), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(new_n809), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1022), .A2(new_n1018), .A3(new_n793), .A4(new_n1024), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT123), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1088), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1142), .A2(KEYINPUT124), .B1(new_n1088), .B2(G168), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1141), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1140), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1145));
  OAI21_X1  g720(.A(G8), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT51), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G168), .A2(new_n1088), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT51), .B(new_n1150), .C1(new_n1138), .C2(G8), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1150), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1135), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1085), .A2(new_n1087), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G288), .A2(G1976), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1106), .A2(new_n1157), .B1(new_n1097), .B2(new_n592), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1089), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1107), .A2(new_n1113), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT113), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1108), .A2(new_n1161), .A3(new_n1116), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1111), .B1(G8), .B2(new_n1112), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT113), .B1(new_n1163), .B2(new_n1107), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1088), .B(G286), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1113), .A2(new_n1165), .A3(KEYINPUT63), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1108), .A2(new_n1165), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1160), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1150), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1142), .A2(KEYINPUT124), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1151), .B1(new_n1176), .B2(KEYINPUT51), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1154), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT62), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1153), .A2(new_n1180), .A3(new_n1154), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1117), .A2(G171), .A3(new_n1131), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1156), .A2(new_n1173), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n755), .B(new_n762), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n820), .B(G1996), .ZN(new_n1188));
  INV_X1    g763(.A(new_n738), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n736), .A2(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n736), .A2(new_n1189), .ZN(new_n1191));
  NOR4_X1   g766(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(G1986), .B2(G290), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n604), .A2(new_n727), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1185), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1184), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT48), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1193), .B2(new_n1185), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1054), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT46), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1185), .B1(new_n1187), .B2(new_n820), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT47), .Z(new_n1203));
  NAND4_X1  g778(.A1(new_n1192), .A2(new_n1197), .A3(new_n727), .A4(new_n604), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1190), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1204), .B(new_n1206), .C1(G2067), .C2(new_n755), .ZN(new_n1207));
  AOI211_X1 g782(.A(new_n1198), .B(new_n1203), .C1(new_n1185), .C2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1196), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g784(.A(G319), .ZN(new_n1211));
  NOR3_X1   g785(.A1(G401), .A2(new_n1211), .A3(G227), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n705), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n1213), .B1(new_n895), .B2(new_n898), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n998), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1216));
  AND3_X1   g790(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1215), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1217), .A2(new_n1218), .ZN(G308));
  NAND2_X1  g793(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n1220), .A2(KEYINPUT127), .ZN(new_n1221));
  NAND3_X1  g795(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1222), .ZN(G225));
endmodule


