

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G651), .A2(n582), .ZN(n786) );
  XNOR2_X1 U554 ( .A(n534), .B(n533), .ZN(G164) );
  NOR2_X4 U555 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X1 U556 ( .A(n525), .B(n524), .ZN(n536) );
  AND2_X1 U557 ( .A1(n536), .A2(G138), .ZN(n527) );
  NOR2_X1 U558 ( .A1(n719), .A2(n734), .ZN(n521) );
  AND2_X1 U559 ( .A1(n679), .A2(G1996), .ZN(n635) );
  NOR2_X1 U560 ( .A1(n648), .A2(n1001), .ZN(n664) );
  INV_X1 U561 ( .A(KEYINPUT97), .ZN(n693) );
  INV_X1 U562 ( .A(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n603) );
  XNOR2_X1 U564 ( .A(n603), .B(KEYINPUT64), .ZN(n632) );
  INV_X1 U565 ( .A(KEYINPUT89), .ZN(n526) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n789) );
  INV_X1 U567 ( .A(G2105), .ZN(n530) );
  AND2_X1 U568 ( .A1(n530), .A2(G2104), .ZN(n867) );
  NAND2_X1 U569 ( .A1(G102), .A2(n867), .ZN(n523) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n870) );
  NAND2_X1 U571 ( .A1(G114), .A2(n870), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n529) );
  XNOR2_X1 U573 ( .A(n527), .B(n526), .ZN(n528) );
  NOR2_X1 U574 ( .A1(n529), .A2(n528), .ZN(n532) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n530), .ZN(n871) );
  NAND2_X1 U576 ( .A1(n871), .A2(G126), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n532), .A2(n531), .ZN(n534) );
  INV_X1 U578 ( .A(KEYINPUT90), .ZN(n533) );
  NAND2_X1 U579 ( .A1(G101), .A2(n867), .ZN(n535) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n535), .Z(n540) );
  INV_X1 U581 ( .A(n536), .ZN(n537) );
  INV_X1 U582 ( .A(n537), .ZN(n866) );
  NAND2_X1 U583 ( .A1(n866), .A2(G137), .ZN(n538) );
  XOR2_X1 U584 ( .A(KEYINPUT65), .B(n538), .Z(n539) );
  NAND2_X1 U585 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U586 ( .A1(G113), .A2(n870), .ZN(n542) );
  NAND2_X1 U587 ( .A1(G125), .A2(n871), .ZN(n541) );
  NAND2_X1 U588 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U589 ( .A1(n544), .A2(n543), .ZN(G160) );
  NAND2_X1 U590 ( .A1(G89), .A2(n789), .ZN(n545) );
  XNOR2_X1 U591 ( .A(n545), .B(KEYINPUT4), .ZN(n546) );
  XNOR2_X1 U592 ( .A(n546), .B(KEYINPUT76), .ZN(n548) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n582) );
  INV_X1 U594 ( .A(G651), .ZN(n551) );
  NOR2_X1 U595 ( .A1(n582), .A2(n551), .ZN(n790) );
  NAND2_X1 U596 ( .A1(G76), .A2(n790), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U598 ( .A(n549), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U599 ( .A1(n786), .A2(G51), .ZN(n550) );
  XOR2_X1 U600 ( .A(KEYINPUT77), .B(n550), .Z(n554) );
  NOR2_X1 U601 ( .A1(G543), .A2(n551), .ZN(n552) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n552), .Z(n785) );
  NAND2_X1 U603 ( .A1(n785), .A2(G63), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U606 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U607 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G91), .A2(n789), .ZN(n560) );
  NAND2_X1 U610 ( .A1(G78), .A2(n790), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U612 ( .A(KEYINPUT66), .B(n561), .Z(n567) );
  NAND2_X1 U613 ( .A1(n786), .A2(G53), .ZN(n562) );
  XOR2_X1 U614 ( .A(KEYINPUT67), .B(n562), .Z(n564) );
  NAND2_X1 U615 ( .A1(n785), .A2(G65), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U617 ( .A(KEYINPUT68), .B(n565), .Z(n566) );
  NAND2_X1 U618 ( .A1(n567), .A2(n566), .ZN(G299) );
  NAND2_X1 U619 ( .A1(G64), .A2(n785), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G52), .A2(n786), .ZN(n568) );
  NAND2_X1 U621 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U622 ( .A1(G90), .A2(n789), .ZN(n571) );
  NAND2_X1 U623 ( .A1(G77), .A2(n790), .ZN(n570) );
  NAND2_X1 U624 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n572), .Z(n573) );
  NOR2_X1 U626 ( .A1(n574), .A2(n573), .ZN(G171) );
  NAND2_X1 U627 ( .A1(G62), .A2(n785), .ZN(n576) );
  NAND2_X1 U628 ( .A1(G50), .A2(n786), .ZN(n575) );
  NAND2_X1 U629 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U630 ( .A(KEYINPUT86), .B(n577), .Z(n581) );
  NAND2_X1 U631 ( .A1(G88), .A2(n789), .ZN(n579) );
  NAND2_X1 U632 ( .A1(G75), .A2(n790), .ZN(n578) );
  AND2_X1 U633 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n581), .A2(n580), .ZN(G303) );
  NAND2_X1 U635 ( .A1(G87), .A2(n582), .ZN(n583) );
  XNOR2_X1 U636 ( .A(n583), .B(KEYINPUT84), .ZN(n588) );
  NAND2_X1 U637 ( .A1(G49), .A2(n786), .ZN(n585) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n785), .A2(n586), .ZN(n587) );
  NAND2_X1 U641 ( .A1(n588), .A2(n587), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G73), .A2(n790), .ZN(n589) );
  XNOR2_X1 U643 ( .A(n589), .B(KEYINPUT2), .ZN(n596) );
  NAND2_X1 U644 ( .A1(G61), .A2(n785), .ZN(n591) );
  NAND2_X1 U645 ( .A1(G48), .A2(n786), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U647 ( .A1(G86), .A2(n789), .ZN(n592) );
  XNOR2_X1 U648 ( .A(KEYINPUT85), .B(n592), .ZN(n593) );
  NOR2_X1 U649 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U650 ( .A1(n596), .A2(n595), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G85), .A2(n789), .ZN(n598) );
  NAND2_X1 U652 ( .A1(G72), .A2(n790), .ZN(n597) );
  NAND2_X1 U653 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U654 ( .A1(G60), .A2(n785), .ZN(n600) );
  NAND2_X1 U655 ( .A1(G47), .A2(n786), .ZN(n599) );
  NAND2_X1 U656 ( .A1(n600), .A2(n599), .ZN(n601) );
  OR2_X1 U657 ( .A1(n602), .A2(n601), .ZN(G290) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n634) );
  NOR2_X1 U659 ( .A1(n634), .A2(n632), .ZN(n753) );
  XNOR2_X1 U660 ( .A(G2067), .B(KEYINPUT37), .ZN(n751) );
  NAND2_X1 U661 ( .A1(G140), .A2(n866), .ZN(n605) );
  NAND2_X1 U662 ( .A1(G104), .A2(n867), .ZN(n604) );
  NAND2_X1 U663 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U664 ( .A(KEYINPUT34), .B(n606), .ZN(n611) );
  NAND2_X1 U665 ( .A1(G116), .A2(n870), .ZN(n608) );
  NAND2_X1 U666 ( .A1(G128), .A2(n871), .ZN(n607) );
  NAND2_X1 U667 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U668 ( .A(KEYINPUT35), .B(n609), .Z(n610) );
  NOR2_X1 U669 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U670 ( .A(KEYINPUT36), .B(n612), .ZN(n878) );
  NOR2_X1 U671 ( .A1(n751), .A2(n878), .ZN(n974) );
  NAND2_X1 U672 ( .A1(n753), .A2(n974), .ZN(n749) );
  NAND2_X1 U673 ( .A1(G107), .A2(n870), .ZN(n614) );
  NAND2_X1 U674 ( .A1(G119), .A2(n871), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U676 ( .A(KEYINPUT91), .B(n615), .ZN(n619) );
  NAND2_X1 U677 ( .A1(n866), .A2(G131), .ZN(n617) );
  NAND2_X1 U678 ( .A1(G95), .A2(n867), .ZN(n616) );
  AND2_X1 U679 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U680 ( .A1(n619), .A2(n618), .ZN(n880) );
  NAND2_X1 U681 ( .A1(G1991), .A2(n880), .ZN(n629) );
  NAND2_X1 U682 ( .A1(G105), .A2(n867), .ZN(n620) );
  XNOR2_X1 U683 ( .A(n620), .B(KEYINPUT38), .ZN(n627) );
  NAND2_X1 U684 ( .A1(G141), .A2(n866), .ZN(n622) );
  NAND2_X1 U685 ( .A1(G117), .A2(n870), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U687 ( .A1(n871), .A2(G129), .ZN(n623) );
  XOR2_X1 U688 ( .A(KEYINPUT92), .B(n623), .Z(n624) );
  NOR2_X1 U689 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U690 ( .A1(n627), .A2(n626), .ZN(n879) );
  NAND2_X1 U691 ( .A1(G1996), .A2(n879), .ZN(n628) );
  NAND2_X1 U692 ( .A1(n629), .A2(n628), .ZN(n967) );
  NAND2_X1 U693 ( .A1(n967), .A2(n753), .ZN(n630) );
  XNOR2_X1 U694 ( .A(n630), .B(KEYINPUT93), .ZN(n746) );
  INV_X1 U695 ( .A(n746), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n749), .A2(n631), .ZN(n741) );
  INV_X1 U697 ( .A(n632), .ZN(n633) );
  NOR2_X4 U698 ( .A1(n634), .A2(n633), .ZN(n679) );
  XOR2_X1 U699 ( .A(KEYINPUT26), .B(n635), .Z(n637) );
  INV_X1 U700 ( .A(n679), .ZN(n695) );
  NAND2_X1 U701 ( .A1(n695), .A2(G1341), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n637), .A2(n636), .ZN(n648) );
  NAND2_X1 U703 ( .A1(n789), .A2(G81), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n638), .B(KEYINPUT12), .ZN(n640) );
  NAND2_X1 U705 ( .A1(G68), .A2(n790), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U707 ( .A(KEYINPUT13), .B(n641), .Z(n645) );
  NAND2_X1 U708 ( .A1(G56), .A2(n785), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT71), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n643), .B(KEYINPUT14), .ZN(n644) );
  NOR2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U712 ( .A1(n786), .A2(G43), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n1001) );
  NAND2_X1 U714 ( .A1(G79), .A2(n790), .ZN(n650) );
  NAND2_X1 U715 ( .A1(G54), .A2(n786), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT73), .ZN(n653) );
  NAND2_X1 U718 ( .A1(G66), .A2(n785), .ZN(n652) );
  NAND2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U720 ( .A1(n789), .A2(G92), .ZN(n654) );
  XOR2_X1 U721 ( .A(KEYINPUT72), .B(n654), .Z(n655) );
  NOR2_X1 U722 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U723 ( .A(n657), .B(KEYINPUT15), .Z(n658) );
  XNOR2_X1 U724 ( .A(KEYINPUT74), .B(n658), .ZN(n1000) );
  NAND2_X1 U725 ( .A1(n664), .A2(n1000), .ZN(n663) );
  INV_X1 U726 ( .A(G2067), .ZN(n945) );
  NOR2_X1 U727 ( .A1(n695), .A2(n945), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n659), .B(KEYINPUT95), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n695), .A2(G1348), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n666) );
  OR2_X1 U732 ( .A1(n1000), .A2(n664), .ZN(n665) );
  NAND2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT96), .ZN(n672) );
  NAND2_X1 U735 ( .A1(n679), .A2(G2072), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n668), .B(KEYINPUT27), .ZN(n670) );
  INV_X1 U737 ( .A(G1956), .ZN(n927) );
  NOR2_X1 U738 ( .A1(n927), .A2(n679), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n673) );
  INV_X1 U740 ( .A(G299), .ZN(n1008) );
  NAND2_X1 U741 ( .A1(n673), .A2(n1008), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n673), .A2(n1008), .ZN(n674) );
  XOR2_X1 U744 ( .A(n674), .B(KEYINPUT28), .Z(n675) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U746 ( .A(KEYINPUT29), .B(n677), .Z(n683) );
  OR2_X1 U747 ( .A1(n679), .A2(G1961), .ZN(n681) );
  XNOR2_X1 U748 ( .A(G2078), .B(KEYINPUT25), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n678), .B(KEYINPUT94), .ZN(n952) );
  NAND2_X1 U750 ( .A1(n679), .A2(n952), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n687), .A2(G171), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n692) );
  NAND2_X1 U754 ( .A1(G8), .A2(n695), .ZN(n734) );
  NOR2_X1 U755 ( .A1(G1966), .A2(n734), .ZN(n708) );
  NOR2_X1 U756 ( .A1(G2084), .A2(n695), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n708), .A2(n705), .ZN(n684) );
  NAND2_X1 U758 ( .A1(G8), .A2(n684), .ZN(n685) );
  XNOR2_X1 U759 ( .A(KEYINPUT30), .B(n685), .ZN(n686) );
  NOR2_X1 U760 ( .A1(G168), .A2(n686), .ZN(n689) );
  NOR2_X1 U761 ( .A1(G171), .A2(n687), .ZN(n688) );
  NOR2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U763 ( .A(KEYINPUT31), .B(n690), .Z(n691) );
  NAND2_X1 U764 ( .A1(n692), .A2(n691), .ZN(n706) );
  NAND2_X1 U765 ( .A1(G286), .A2(n706), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n694), .B(n693), .ZN(n701) );
  NOR2_X1 U767 ( .A1(G2090), .A2(n695), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n696), .B(KEYINPUT98), .ZN(n698) );
  NOR2_X1 U769 ( .A1(n734), .A2(G1971), .ZN(n697) );
  NOR2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U771 ( .A1(G303), .A2(n699), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n702), .A2(G8), .ZN(n704) );
  XOR2_X1 U774 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n703) );
  XNOR2_X1 U775 ( .A(n704), .B(n703), .ZN(n712) );
  NAND2_X1 U776 ( .A1(G8), .A2(n705), .ZN(n710) );
  INV_X1 U777 ( .A(n706), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n733) );
  NOR2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  NOR2_X1 U782 ( .A1(G1971), .A2(G303), .ZN(n713) );
  XNOR2_X1 U783 ( .A(KEYINPUT100), .B(n713), .ZN(n714) );
  NOR2_X1 U784 ( .A1(n1013), .A2(n714), .ZN(n716) );
  INV_X1 U785 ( .A(KEYINPUT33), .ZN(n715) );
  AND2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n733), .A2(n717), .ZN(n725) );
  NAND2_X1 U788 ( .A1(G288), .A2(G1976), .ZN(n718) );
  XOR2_X1 U789 ( .A(KEYINPUT101), .B(n718), .Z(n1006) );
  INV_X1 U790 ( .A(n1006), .ZN(n719) );
  NOR2_X1 U791 ( .A1(KEYINPUT33), .A2(n521), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n1013), .A2(KEYINPUT33), .ZN(n720) );
  NOR2_X1 U793 ( .A1(n720), .A2(n734), .ZN(n721) );
  NOR2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U795 ( .A(G1981), .B(G305), .Z(n997) );
  AND2_X1 U796 ( .A1(n723), .A2(n997), .ZN(n724) );
  AND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n739) );
  NOR2_X1 U798 ( .A1(G2090), .A2(G303), .ZN(n726) );
  NAND2_X1 U799 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U800 ( .A(n727), .B(KEYINPUT102), .ZN(n731) );
  NOR2_X1 U801 ( .A1(G1981), .A2(G305), .ZN(n728) );
  XOR2_X1 U802 ( .A(n728), .B(KEYINPUT24), .Z(n729) );
  NOR2_X1 U803 ( .A1(n734), .A2(n729), .ZN(n735) );
  INV_X1 U804 ( .A(n735), .ZN(n730) );
  AND2_X1 U805 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n737) );
  OR2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n1012) );
  NAND2_X1 U812 ( .A1(n1012), .A2(n753), .ZN(n742) );
  NAND2_X1 U813 ( .A1(n743), .A2(n742), .ZN(n756) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n879), .ZN(n977) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n880), .ZN(n968) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n744) );
  NOR2_X1 U817 ( .A1(n968), .A2(n744), .ZN(n745) );
  NOR2_X1 U818 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U819 ( .A1(n977), .A2(n747), .ZN(n748) );
  XNOR2_X1 U820 ( .A(n748), .B(KEYINPUT39), .ZN(n750) );
  NAND2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U822 ( .A1(n751), .A2(n878), .ZN(n982) );
  NAND2_X1 U823 ( .A1(n752), .A2(n982), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U825 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U826 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U828 ( .A(G57), .ZN(G237) );
  INV_X1 U829 ( .A(G82), .ZN(G220) );
  NAND2_X1 U830 ( .A1(G7), .A2(G661), .ZN(n758) );
  XNOR2_X1 U831 ( .A(n758), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U832 ( .A(G223), .B(KEYINPUT70), .Z(n819) );
  NAND2_X1 U833 ( .A1(n819), .A2(G567), .ZN(n759) );
  XOR2_X1 U834 ( .A(KEYINPUT11), .B(n759), .Z(G234) );
  INV_X1 U835 ( .A(G860), .ZN(n827) );
  OR2_X1 U836 ( .A1(n1001), .A2(n827), .ZN(G153) );
  NOR2_X1 U837 ( .A1(G868), .A2(n1000), .ZN(n761) );
  INV_X1 U838 ( .A(G868), .ZN(n802) );
  NOR2_X1 U839 ( .A1(G171), .A2(n802), .ZN(n760) );
  NOR2_X1 U840 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U841 ( .A(KEYINPUT75), .B(n762), .ZN(G284) );
  XNOR2_X1 U842 ( .A(KEYINPUT78), .B(n802), .ZN(n763) );
  NOR2_X1 U843 ( .A1(G286), .A2(n763), .ZN(n765) );
  NOR2_X1 U844 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U845 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U846 ( .A1(n827), .A2(G559), .ZN(n766) );
  NAND2_X1 U847 ( .A1(n766), .A2(n1000), .ZN(n767) );
  XNOR2_X1 U848 ( .A(n767), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U849 ( .A1(G868), .A2(n1001), .ZN(n768) );
  XOR2_X1 U850 ( .A(KEYINPUT79), .B(n768), .Z(n772) );
  NAND2_X1 U851 ( .A1(G868), .A2(n1000), .ZN(n769) );
  NOR2_X1 U852 ( .A1(G559), .A2(n769), .ZN(n770) );
  XNOR2_X1 U853 ( .A(KEYINPUT80), .B(n770), .ZN(n771) );
  NOR2_X1 U854 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U855 ( .A1(G99), .A2(n867), .ZN(n774) );
  NAND2_X1 U856 ( .A1(G111), .A2(n870), .ZN(n773) );
  NAND2_X1 U857 ( .A1(n774), .A2(n773), .ZN(n781) );
  NAND2_X1 U858 ( .A1(n866), .A2(G135), .ZN(n775) );
  XNOR2_X1 U859 ( .A(KEYINPUT81), .B(n775), .ZN(n778) );
  NAND2_X1 U860 ( .A1(n871), .A2(G123), .ZN(n776) );
  XOR2_X1 U861 ( .A(KEYINPUT18), .B(n776), .Z(n777) );
  NOR2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U863 ( .A(KEYINPUT82), .B(n779), .Z(n780) );
  NOR2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n970) );
  XNOR2_X1 U865 ( .A(G2096), .B(n970), .ZN(n783) );
  INV_X1 U866 ( .A(G2100), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(G156) );
  INV_X1 U868 ( .A(G303), .ZN(G166) );
  NAND2_X1 U869 ( .A1(n1000), .A2(G559), .ZN(n784) );
  XOR2_X1 U870 ( .A(n1001), .B(n784), .Z(n826) );
  XNOR2_X1 U871 ( .A(n1008), .B(G166), .ZN(n800) );
  XNOR2_X1 U872 ( .A(KEYINPUT19), .B(G288), .ZN(n796) );
  NAND2_X1 U873 ( .A1(G67), .A2(n785), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G55), .A2(n786), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n794) );
  NAND2_X1 U876 ( .A1(G93), .A2(n789), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G80), .A2(n790), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U880 ( .A(n795), .B(KEYINPUT83), .ZN(n828) );
  XNOR2_X1 U881 ( .A(n796), .B(n828), .ZN(n797) );
  XNOR2_X1 U882 ( .A(n797), .B(G290), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n798), .B(G305), .ZN(n799) );
  XNOR2_X1 U884 ( .A(n800), .B(n799), .ZN(n894) );
  XNOR2_X1 U885 ( .A(n826), .B(n894), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n801), .A2(G868), .ZN(n804) );
  NAND2_X1 U887 ( .A1(n802), .A2(n828), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2084), .A2(G2078), .ZN(n805) );
  XNOR2_X1 U890 ( .A(n805), .B(KEYINPUT87), .ZN(n806) );
  XNOR2_X1 U891 ( .A(KEYINPUT20), .B(n806), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n807), .A2(G2090), .ZN(n808) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(n808), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n809), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U896 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NAND2_X1 U897 ( .A1(G483), .A2(G661), .ZN(n817) );
  NOR2_X1 U898 ( .A1(G220), .A2(G219), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT22), .B(n810), .Z(n811) );
  NOR2_X1 U900 ( .A1(G218), .A2(n811), .ZN(n812) );
  NAND2_X1 U901 ( .A1(G96), .A2(n812), .ZN(n824) );
  NAND2_X1 U902 ( .A1(n824), .A2(G2106), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G69), .A2(G120), .ZN(n813) );
  NOR2_X1 U904 ( .A1(G237), .A2(n813), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G108), .A2(n814), .ZN(n825) );
  NAND2_X1 U906 ( .A1(n825), .A2(G567), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n849) );
  NOR2_X1 U908 ( .A1(n817), .A2(n849), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n818), .B(KEYINPUT88), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G36), .A2(n823), .ZN(G176) );
  NAND2_X1 U911 ( .A1(n819), .A2(G2106), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n820), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U914 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(G188) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(n828), .ZN(G145) );
  XOR2_X1 U925 ( .A(KEYINPUT105), .B(G2090), .Z(n831) );
  XNOR2_X1 U926 ( .A(G2078), .B(G2072), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U928 ( .A(n832), .B(G2096), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2084), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U931 ( .A(KEYINPUT43), .B(G2678), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2100), .B(KEYINPUT42), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(n838), .B(n837), .Z(G227) );
  XNOR2_X1 U935 ( .A(G1996), .B(KEYINPUT106), .ZN(n848) );
  XOR2_X1 U936 ( .A(G1981), .B(G1956), .Z(n840) );
  XNOR2_X1 U937 ( .A(G1991), .B(G1961), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2474), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(G229) );
  INV_X1 U946 ( .A(n849), .ZN(G319) );
  NAND2_X1 U947 ( .A1(G124), .A2(n871), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G100), .A2(n867), .ZN(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT107), .B(n851), .Z(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G136), .A2(n866), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G112), .A2(n870), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U955 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U956 ( .A1(G118), .A2(n870), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G130), .A2(n871), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U959 ( .A1(n867), .A2(G106), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT108), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G142), .A2(n866), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U963 ( .A(KEYINPUT45), .B(n863), .Z(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n890) );
  NAND2_X1 U965 ( .A1(G139), .A2(n866), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G103), .A2(n867), .ZN(n868) );
  NAND2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U968 ( .A1(G115), .A2(n870), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G127), .A2(n871), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n984) );
  XOR2_X1 U973 ( .A(G160), .B(n984), .Z(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(n883) );
  XNOR2_X1 U975 ( .A(G162), .B(n879), .ZN(n881) );
  XNOR2_X1 U976 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U977 ( .A(n883), .B(n882), .Z(n888) );
  XOR2_X1 U978 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U979 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U981 ( .A(KEYINPUT48), .B(n886), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U983 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U984 ( .A(G164), .B(n891), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n892), .B(n970), .ZN(n893) );
  NOR2_X1 U986 ( .A1(G37), .A2(n893), .ZN(G395) );
  INV_X1 U987 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U988 ( .A(n1001), .B(n894), .ZN(n896) );
  XNOR2_X1 U989 ( .A(G301), .B(n1000), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U991 ( .A(G286), .B(n897), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G397) );
  XNOR2_X1 U993 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n912) );
  XOR2_X1 U996 ( .A(KEYINPUT103), .B(G2427), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2435), .B(G2438), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n909) );
  XOR2_X1 U999 ( .A(G2443), .B(G2430), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G2454), .B(G2446), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1002 ( .A(n905), .B(G2451), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n910), .A2(G14), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n915), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1014 ( .A(KEYINPUT123), .B(G16), .ZN(n941) );
  XNOR2_X1 U1015 ( .A(G1971), .B(G22), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G23), .B(G1976), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n919) );
  XOR2_X1 U1018 ( .A(G1986), .B(G24), .Z(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G21), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G1961), .B(G5), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n938) );
  XNOR2_X1 U1026 ( .A(KEYINPUT59), .B(G1348), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n926), .B(G4), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(G20), .B(n927), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G1341), .B(G19), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G1981), .B(G6), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1033 ( .A(KEYINPUT124), .B(n932), .Z(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1035 ( .A(KEYINPUT125), .B(n935), .Z(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT60), .B(n936), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(KEYINPUT61), .B(n939), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n1027) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(KEYINPUT55), .ZN(n962) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n942) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n942), .ZN(n959) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1044 ( .A(G1996), .B(G32), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G26), .B(n945), .ZN(n946) );
  NAND2_X1 U1048 ( .A1(n946), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1049 ( .A(G25), .B(G1991), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(KEYINPUT116), .B(n947), .ZN(n948) );
  NOR2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1053 ( .A(n952), .B(G27), .Z(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n960), .B(KEYINPUT118), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1060 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n965), .A2(G11), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n966), .B(KEYINPUT119), .ZN(n996) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G2084), .B(G160), .Z(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(KEYINPUT113), .B(n975), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT51), .B(n978), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n981), .B(KEYINPUT114), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(G2072), .B(n984), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G164), .B(G2078), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT50), .B(n987), .Z(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT115), .B(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT52), .B(n991), .ZN(n993) );
  INV_X1 U1083 ( .A(KEYINPUT55), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(G29), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1025) );
  XNOR2_X1 U1087 ( .A(KEYINPUT56), .B(G16), .ZN(n1022) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G168), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(n999), .B(KEYINPUT57), .ZN(n1020) );
  XNOR2_X1 U1091 ( .A(G1348), .B(n1000), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G301), .B(G1961), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1001), .B(G1341), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1018) );
  XNOR2_X1 U1096 ( .A(G166), .B(G1971), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(G1956), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT120), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT121), .B(n1016), .Z(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT122), .B(n1023), .Z(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

