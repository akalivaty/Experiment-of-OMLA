

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746;

  NAND2_X1 U366 ( .A1(n630), .A2(n629), .ZN(n633) );
  NOR2_X1 U367 ( .A1(G953), .A2(G237), .ZN(n528) );
  XOR2_X1 U368 ( .A(n501), .B(KEYINPUT24), .Z(n346) );
  XNOR2_X2 U369 ( .A(n360), .B(n390), .ZN(n369) );
  NOR2_X2 U370 ( .A1(n701), .A2(G902), .ZN(n464) );
  XNOR2_X2 U371 ( .A(n487), .B(G137), .ZN(n488) );
  XNOR2_X2 U372 ( .A(n500), .B(n489), .ZN(n728) );
  NOR2_X1 U373 ( .A1(n419), .A2(n721), .ZN(n655) );
  NAND2_X1 U374 ( .A1(n365), .A2(n362), .ZN(n420) );
  AND2_X1 U375 ( .A1(n367), .A2(n353), .ZN(n365) );
  NAND2_X1 U376 ( .A1(n364), .A2(n363), .ZN(n362) );
  NAND2_X1 U377 ( .A1(n391), .A2(n352), .ZN(n360) );
  AND2_X2 U378 ( .A1(n658), .A2(n352), .ZN(n712) );
  XNOR2_X1 U379 ( .A(n373), .B(n583), .ZN(n617) );
  NOR2_X1 U380 ( .A1(n436), .A2(n434), .ZN(n443) );
  XNOR2_X1 U381 ( .A(n375), .B(KEYINPUT0), .ZN(n605) );
  NOR2_X1 U382 ( .A1(n582), .A2(n581), .ZN(n375) );
  XNOR2_X1 U383 ( .A(n603), .B(n542), .ZN(n601) );
  XNOR2_X1 U384 ( .A(n506), .B(KEYINPUT20), .ZN(n511) );
  XNOR2_X1 U385 ( .A(n515), .B(n514), .ZN(n518) );
  XNOR2_X1 U386 ( .A(n407), .B(G119), .ZN(n527) );
  XNOR2_X1 U387 ( .A(n415), .B(G104), .ZN(n372) );
  XNOR2_X1 U388 ( .A(KEYINPUT4), .B(KEYINPUT70), .ZN(n486) );
  XOR2_X1 U389 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n515) );
  NOR2_X1 U390 ( .A1(n419), .A2(n721), .ZN(n347) );
  XNOR2_X1 U391 ( .A(n397), .B(n433), .ZN(n431) );
  XNOR2_X1 U392 ( .A(n534), .B(n447), .ZN(n695) );
  AND2_X1 U393 ( .A1(n430), .A2(KEYINPUT75), .ZN(n423) );
  XNOR2_X1 U394 ( .A(n729), .B(G146), .ZN(n534) );
  XOR2_X1 U395 ( .A(G101), .B(G110), .Z(n492) );
  XNOR2_X1 U396 ( .A(n409), .B(G116), .ZN(n483) );
  XNOR2_X1 U397 ( .A(G122), .B(G107), .ZN(n409) );
  XNOR2_X1 U398 ( .A(n484), .B(n724), .ZN(n660) );
  INV_X1 U399 ( .A(KEYINPUT84), .ZN(n433) );
  NAND2_X1 U400 ( .A1(n746), .A2(n560), .ZN(n397) );
  AND2_X1 U401 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U402 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U403 ( .A1(n421), .A2(KEYINPUT71), .ZN(n382) );
  INV_X1 U404 ( .A(n617), .ZN(n628) );
  XNOR2_X1 U405 ( .A(G125), .B(G146), .ZN(n478) );
  XNOR2_X1 U406 ( .A(n402), .B(n401), .ZN(n498) );
  INV_X1 U407 ( .A(KEYINPUT8), .ZN(n401) );
  NAND2_X1 U408 ( .A1(n450), .A2(n448), .ZN(n616) );
  NOR2_X1 U409 ( .A1(n692), .A2(n449), .ZN(n448) );
  XNOR2_X1 U410 ( .A(n386), .B(n451), .ZN(n450) );
  INV_X1 U411 ( .A(n694), .ZN(n449) );
  XNOR2_X1 U412 ( .A(G107), .B(G104), .ZN(n491) );
  NAND2_X1 U413 ( .A1(n435), .A2(n348), .ZN(n434) );
  NAND2_X1 U414 ( .A1(n633), .A2(n513), .ZN(n437) );
  INV_X1 U415 ( .A(KEYINPUT30), .ZN(n441) );
  XNOR2_X1 U416 ( .A(n527), .B(n406), .ZN(n530) );
  INV_X1 U417 ( .A(KEYINPUT96), .ZN(n406) );
  XNOR2_X1 U418 ( .A(G128), .B(G140), .ZN(n501) );
  XNOR2_X1 U419 ( .A(n478), .B(KEYINPUT10), .ZN(n500) );
  XNOR2_X1 U420 ( .A(n503), .B(n502), .ZN(n395) );
  XOR2_X1 U421 ( .A(KEYINPUT23), .B(G137), .Z(n503) );
  BUF_X1 U422 ( .A(n595), .Z(n408) );
  NAND2_X1 U423 ( .A1(n601), .A2(n370), .ZN(n571) );
  NOR2_X1 U424 ( .A1(n371), .A2(n568), .ZN(n370) );
  INV_X1 U425 ( .A(KEYINPUT102), .ZN(n473) );
  NOR2_X1 U426 ( .A1(n571), .A2(n546), .ZN(n400) );
  INV_X1 U427 ( .A(KEYINPUT36), .ZN(n399) );
  INV_X1 U428 ( .A(n601), .ZN(n591) );
  OR2_X1 U429 ( .A1(n589), .A2(n630), .ZN(n403) );
  XNOR2_X1 U430 ( .A(n417), .B(n355), .ZN(n594) );
  NOR2_X1 U431 ( .A1(n622), .A2(n541), .ZN(n418) );
  XNOR2_X1 U432 ( .A(n454), .B(G475), .ZN(n453) );
  INV_X1 U433 ( .A(KEYINPUT13), .ZN(n454) );
  XNOR2_X1 U434 ( .A(n472), .B(n349), .ZN(n540) );
  NOR2_X1 U435 ( .A1(G902), .A2(n710), .ZN(n472) );
  XNOR2_X1 U436 ( .A(n605), .B(n374), .ZN(n608) );
  INV_X1 U437 ( .A(KEYINPUT93), .ZN(n374) );
  INV_X1 U438 ( .A(G472), .ZN(n396) );
  XNOR2_X1 U439 ( .A(n412), .B(n482), .ZN(n724) );
  XNOR2_X1 U440 ( .A(n413), .B(n483), .ZN(n412) );
  XNOR2_X1 U441 ( .A(n372), .B(n414), .ZN(n413) );
  INV_X1 U442 ( .A(n408), .ZN(n632) );
  NAND2_X1 U443 ( .A1(n426), .A2(n428), .ZN(n425) );
  INV_X1 U444 ( .A(KEYINPUT75), .ZN(n428) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n514) );
  NAND2_X1 U446 ( .A1(n389), .A2(n387), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n388), .B(n356), .ZN(n387) );
  NAND2_X1 U448 ( .A1(n383), .A2(n380), .ZN(n389) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n451) );
  XNOR2_X1 U450 ( .A(G143), .B(KEYINPUT12), .ZN(n458) );
  XOR2_X1 U451 ( .A(KEYINPUT4), .B(KEYINPUT70), .Z(n475) );
  XNOR2_X1 U452 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n476) );
  OR2_X1 U453 ( .A1(G902), .A2(G237), .ZN(n536) );
  XNOR2_X1 U454 ( .A(n394), .B(n446), .ZN(n595) );
  INV_X1 U455 ( .A(KEYINPUT1), .ZN(n446) );
  NOR2_X1 U456 ( .A1(n604), .A2(n591), .ZN(n373) );
  XNOR2_X1 U457 ( .A(n444), .B(KEYINPUT78), .ZN(n604) );
  NAND2_X1 U458 ( .A1(n595), .A2(n445), .ZN(n444) );
  INV_X1 U459 ( .A(n540), .ZN(n564) );
  XOR2_X1 U460 ( .A(KEYINPUT25), .B(KEYINPUT81), .Z(n508) );
  XNOR2_X1 U461 ( .A(G116), .B(G101), .ZN(n521) );
  XOR2_X1 U462 ( .A(G131), .B(G113), .Z(n522) );
  XNOR2_X1 U463 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n523) );
  INV_X1 U464 ( .A(G113), .ZN(n415) );
  INV_X1 U465 ( .A(KEYINPUT16), .ZN(n414) );
  INV_X1 U466 ( .A(KEYINPUT3), .ZN(n407) );
  NOR2_X1 U467 ( .A1(n616), .A2(n392), .ZN(n376) );
  XNOR2_X1 U468 ( .A(n490), .B(n493), .ZN(n447) );
  OR2_X1 U469 ( .A1(n653), .A2(KEYINPUT119), .ZN(n366) );
  XNOR2_X1 U470 ( .A(n537), .B(KEYINPUT80), .ZN(n558) );
  NOR2_X1 U471 ( .A1(n594), .A2(n408), .ZN(n599) );
  XNOR2_X1 U472 ( .A(n395), .B(n346), .ZN(n504) );
  XNOR2_X1 U473 ( .A(n405), .B(n466), .ZN(n710) );
  XOR2_X1 U474 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n465) );
  XNOR2_X1 U475 ( .A(n702), .B(KEYINPUT59), .ZN(n703) );
  XNOR2_X1 U476 ( .A(n660), .B(n659), .ZN(n661) );
  INV_X1 U477 ( .A(KEYINPUT119), .ZN(n363) );
  XNOR2_X1 U478 ( .A(n544), .B(n361), .ZN(n432) );
  INV_X1 U479 ( .A(KEYINPUT110), .ZN(n361) );
  XNOR2_X1 U480 ( .A(n403), .B(KEYINPUT106), .ZN(n590) );
  NAND2_X1 U481 ( .A1(n540), .A2(n563), .ZN(n452) );
  XNOR2_X1 U482 ( .A(n398), .B(KEYINPUT95), .ZN(n610) );
  AND2_X1 U483 ( .A1(n608), .A2(n609), .ZN(n398) );
  XNOR2_X1 U484 ( .A(n416), .B(n350), .ZN(n559) );
  XNOR2_X1 U485 ( .A(KEYINPUT83), .B(n520), .ZN(n348) );
  XOR2_X1 U486 ( .A(KEYINPUT100), .B(G478), .Z(n349) );
  XOR2_X1 U487 ( .A(n485), .B(KEYINPUT82), .Z(n350) );
  INV_X1 U488 ( .A(n633), .ZN(n445) );
  AND2_X1 U489 ( .A1(n553), .A2(n566), .ZN(n351) );
  NAND2_X1 U490 ( .A1(n615), .A2(n376), .ZN(n352) );
  AND2_X1 U491 ( .A1(n366), .A2(n663), .ZN(n353) );
  OR2_X1 U492 ( .A1(n557), .A2(n574), .ZN(n354) );
  XOR2_X1 U493 ( .A(KEYINPUT65), .B(KEYINPUT22), .Z(n355) );
  XOR2_X1 U494 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n356) );
  XNOR2_X1 U495 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n357) );
  XOR2_X1 U496 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n358) );
  XNOR2_X2 U497 ( .A(n359), .B(n510), .ZN(n630) );
  NOR2_X1 U498 ( .A1(n714), .A2(G902), .ZN(n359) );
  XNOR2_X1 U499 ( .A(n432), .B(n357), .ZN(n742) );
  INV_X1 U500 ( .A(n369), .ZN(n364) );
  NAND2_X1 U501 ( .A1(n369), .A2(n368), .ZN(n367) );
  AND2_X1 U502 ( .A1(n653), .A2(KEYINPUT119), .ZN(n368) );
  NAND2_X1 U503 ( .A1(n348), .A2(n547), .ZN(n371) );
  XNOR2_X1 U504 ( .A(n372), .B(n458), .ZN(n462) );
  NAND2_X1 U505 ( .A1(n608), .A2(n617), .ZN(n585) );
  XNOR2_X2 U506 ( .A(n377), .B(KEYINPUT45), .ZN(n615) );
  NAND2_X1 U507 ( .A1(n613), .A2(n614), .ZN(n377) );
  XNOR2_X2 U508 ( .A(n378), .B(KEYINPUT108), .ZN(n746) );
  OR2_X2 U509 ( .A1(n558), .A2(n354), .ZN(n378) );
  XNOR2_X1 U510 ( .A(n467), .B(n379), .ZN(n405) );
  XNOR2_X2 U511 ( .A(n379), .B(n488), .ZN(n729) );
  XNOR2_X2 U512 ( .A(n474), .B(G134), .ZN(n379) );
  INV_X1 U513 ( .A(n424), .ZN(n381) );
  NAND2_X1 U514 ( .A1(n421), .A2(KEYINPUT71), .ZN(n384) );
  NAND2_X1 U515 ( .A1(n424), .A2(KEYINPUT71), .ZN(n385) );
  NAND2_X1 U516 ( .A1(n745), .A2(n744), .ZN(n388) );
  INV_X1 U517 ( .A(KEYINPUT85), .ZN(n390) );
  NAND2_X1 U518 ( .A1(n393), .A2(n392), .ZN(n391) );
  INV_X1 U519 ( .A(KEYINPUT2), .ZN(n392) );
  INV_X1 U520 ( .A(n655), .ZN(n393) );
  NAND2_X1 U521 ( .A1(n663), .A2(G234), .ZN(n402) );
  BUF_X2 U522 ( .A(n552), .Z(n394) );
  XNOR2_X1 U523 ( .A(n400), .B(n399), .ZN(n543) );
  INV_X1 U524 ( .A(n639), .ZN(n603) );
  NAND2_X1 U525 ( .A1(n639), .A2(n620), .ZN(n442) );
  XNOR2_X2 U526 ( .A(n535), .B(n396), .ZN(n639) );
  XNOR2_X1 U527 ( .A(n442), .B(n441), .ZN(n440) );
  NAND2_X1 U528 ( .A1(n439), .A2(n445), .ZN(n438) );
  XNOR2_X2 U529 ( .A(G902), .B(KEYINPUT15), .ZN(n654) );
  NAND2_X1 U530 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X1 U531 ( .A(n505), .B(n504), .ZN(n714) );
  XNOR2_X2 U532 ( .A(n593), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U533 ( .A1(n404), .A2(n351), .ZN(n556) );
  INV_X1 U534 ( .A(n624), .ZN(n404) );
  XNOR2_X2 U535 ( .A(n555), .B(KEYINPUT103), .ZN(n624) );
  NAND2_X1 U536 ( .A1(n429), .A2(n428), .ZN(n427) );
  NOR2_X1 U537 ( .A1(n739), .A2(n597), .ZN(n598) );
  NAND2_X1 U538 ( .A1(n410), .A2(n351), .ZN(n430) );
  XNOR2_X1 U539 ( .A(n561), .B(KEYINPUT76), .ZN(n410) );
  NAND2_X1 U540 ( .A1(n411), .A2(n455), .ZN(n658) );
  NAND2_X1 U541 ( .A1(n347), .A2(n656), .ZN(n411) );
  INV_X1 U542 ( .A(n559), .ZN(n574) );
  NAND2_X1 U543 ( .A1(n559), .A2(n620), .ZN(n546) );
  NAND2_X1 U544 ( .A1(n660), .A2(n654), .ZN(n416) );
  NAND2_X1 U545 ( .A1(n605), .A2(n418), .ZN(n417) );
  XNOR2_X1 U546 ( .A(n419), .B(n732), .ZN(n731) );
  XNOR2_X2 U547 ( .A(n616), .B(KEYINPUT86), .ZN(n419) );
  XNOR2_X1 U548 ( .A(n420), .B(n358), .ZN(G75) );
  NAND2_X1 U549 ( .A1(n422), .A2(n432), .ZN(n421) );
  NAND2_X1 U550 ( .A1(n423), .A2(n431), .ZN(n422) );
  NAND2_X1 U551 ( .A1(n427), .A2(n425), .ZN(n424) );
  INV_X1 U552 ( .A(n430), .ZN(n426) );
  INV_X1 U553 ( .A(n431), .ZN(n429) );
  NOR2_X1 U554 ( .A1(n394), .A2(n633), .ZN(n609) );
  NAND2_X1 U555 ( .A1(n552), .A2(n513), .ZN(n435) );
  NOR2_X1 U556 ( .A1(n552), .A2(n513), .ZN(n439) );
  NAND2_X1 U557 ( .A1(n443), .A2(n440), .ZN(n537) );
  XNOR2_X1 U558 ( .A(n689), .B(n473), .ZN(n554) );
  XNOR2_X1 U559 ( .A(n483), .B(n465), .ZN(n466) );
  XNOR2_X2 U560 ( .A(n452), .B(KEYINPUT101), .ZN(n689) );
  XNOR2_X2 U561 ( .A(n464), .B(n453), .ZN(n563) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n505) );
  NAND2_X2 U563 ( .A1(n471), .A2(n470), .ZN(n474) );
  XOR2_X1 U564 ( .A(n657), .B(KEYINPUT67), .Z(n455) );
  AND2_X1 U565 ( .A1(G224), .A2(n663), .ZN(n456) );
  AND2_X1 U566 ( .A1(G227), .A2(n663), .ZN(n457) );
  XNOR2_X1 U567 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n583) );
  XNOR2_X1 U568 ( .A(n489), .B(n457), .ZN(n490) );
  XNOR2_X1 U569 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U570 ( .A(n456), .B(n479), .ZN(n480) );
  XNOR2_X1 U571 ( .A(n481), .B(n480), .ZN(n484) );
  XNOR2_X1 U572 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U573 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n538) );
  XNOR2_X1 U574 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U575 ( .A(KEYINPUT90), .B(n664), .Z(n705) );
  XOR2_X1 U576 ( .A(G122), .B(KEYINPUT11), .Z(n460) );
  NAND2_X1 U577 ( .A1(n528), .A2(G214), .ZN(n459) );
  XNOR2_X1 U578 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U579 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U580 ( .A(G131), .B(G140), .Z(n489) );
  XNOR2_X1 U581 ( .A(n463), .B(n728), .ZN(n701) );
  INV_X2 U582 ( .A(G953), .ZN(n663) );
  NAND2_X1 U583 ( .A1(G217), .A2(n498), .ZN(n467) );
  INV_X1 U584 ( .A(G128), .ZN(n468) );
  NAND2_X1 U585 ( .A1(n468), .A2(G143), .ZN(n471) );
  INV_X1 U586 ( .A(G143), .ZN(n469) );
  NAND2_X1 U587 ( .A1(n469), .A2(G128), .ZN(n470) );
  XOR2_X1 U588 ( .A(n474), .B(n475), .Z(n477) );
  XNOR2_X1 U589 ( .A(n477), .B(n476), .ZN(n481) );
  INV_X1 U590 ( .A(n478), .ZN(n479) );
  XNOR2_X1 U591 ( .A(n527), .B(n492), .ZN(n482) );
  NAND2_X1 U592 ( .A1(n536), .A2(G210), .ZN(n485) );
  XOR2_X1 U593 ( .A(n574), .B(KEYINPUT38), .Z(n562) );
  INV_X1 U594 ( .A(n486), .ZN(n487) );
  NOR2_X2 U595 ( .A1(G902), .A2(n695), .ZN(n497) );
  XNOR2_X1 U596 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n495) );
  INV_X1 U597 ( .A(G469), .ZN(n494) );
  XNOR2_X2 U598 ( .A(n497), .B(n496), .ZN(n552) );
  NAND2_X1 U599 ( .A1(G221), .A2(n498), .ZN(n499) );
  XNOR2_X1 U600 ( .A(G119), .B(G110), .ZN(n502) );
  NAND2_X1 U601 ( .A1(n654), .A2(G234), .ZN(n506) );
  NAND2_X1 U602 ( .A1(n511), .A2(G217), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U604 ( .A(KEYINPUT94), .B(n509), .ZN(n510) );
  NAND2_X1 U605 ( .A1(n511), .A2(G221), .ZN(n512) );
  XOR2_X1 U606 ( .A(KEYINPUT21), .B(n512), .Z(n629) );
  INV_X1 U607 ( .A(KEYINPUT107), .ZN(n513) );
  NAND2_X1 U608 ( .A1(n518), .A2(G902), .ZN(n516) );
  XNOR2_X1 U609 ( .A(n516), .B(KEYINPUT91), .ZN(n577) );
  NAND2_X1 U610 ( .A1(G953), .A2(n577), .ZN(n517) );
  NOR2_X1 U611 ( .A1(G900), .A2(n517), .ZN(n519) );
  NAND2_X1 U612 ( .A1(n518), .A2(G952), .ZN(n650) );
  NOR2_X1 U613 ( .A1(G953), .A2(n650), .ZN(n576) );
  NOR2_X1 U614 ( .A1(n519), .A2(n576), .ZN(n520) );
  XNOR2_X1 U615 ( .A(n522), .B(n521), .ZN(n526) );
  XOR2_X1 U616 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n524) );
  XNOR2_X1 U617 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n526), .B(n525), .ZN(n532) );
  NAND2_X1 U619 ( .A1(n528), .A2(G210), .ZN(n529) );
  XNOR2_X1 U620 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U622 ( .A(n534), .B(n533), .ZN(n669) );
  NOR2_X1 U623 ( .A1(n669), .A2(G902), .ZN(n535) );
  NAND2_X1 U624 ( .A1(G214), .A2(n536), .ZN(n620) );
  NOR2_X1 U625 ( .A1(n562), .A2(n558), .ZN(n539) );
  XNOR2_X1 U626 ( .A(n539), .B(n538), .ZN(n569) );
  NOR2_X1 U627 ( .A1(n554), .A2(n569), .ZN(n692) );
  XNOR2_X1 U628 ( .A(n408), .B(KEYINPUT89), .ZN(n589) );
  NOR2_X1 U629 ( .A1(n563), .A2(n540), .ZN(n687) );
  INV_X1 U630 ( .A(n687), .ZN(n568) );
  INV_X1 U631 ( .A(n629), .ZN(n541) );
  NOR2_X1 U632 ( .A1(n541), .A2(n630), .ZN(n547) );
  XNOR2_X1 U633 ( .A(KEYINPUT6), .B(KEYINPUT104), .ZN(n542) );
  NOR2_X1 U634 ( .A1(n589), .A2(n543), .ZN(n544) );
  XOR2_X1 U635 ( .A(KEYINPUT19), .B(KEYINPUT68), .Z(n545) );
  XNOR2_X1 U636 ( .A(n546), .B(n545), .ZN(n582) );
  INV_X1 U637 ( .A(n582), .ZN(n553) );
  NAND2_X1 U638 ( .A1(n547), .A2(n348), .ZN(n548) );
  NOR2_X1 U639 ( .A1(n603), .A2(n548), .ZN(n550) );
  XNOR2_X1 U640 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n549) );
  XNOR2_X1 U641 ( .A(n550), .B(n549), .ZN(n551) );
  NOR2_X1 U642 ( .A1(n394), .A2(n551), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n554), .A2(n568), .ZN(n555) );
  NAND2_X1 U644 ( .A1(n556), .A2(KEYINPUT47), .ZN(n560) );
  NOR2_X1 U645 ( .A1(n563), .A2(n564), .ZN(n586) );
  INV_X1 U646 ( .A(n586), .ZN(n557) );
  NOR2_X1 U647 ( .A1(n624), .A2(KEYINPUT47), .ZN(n561) );
  INV_X1 U648 ( .A(n562), .ZN(n619) );
  NAND2_X1 U649 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U650 ( .A1(n564), .A2(n563), .ZN(n622) );
  NOR2_X1 U651 ( .A1(n623), .A2(n622), .ZN(n565) );
  XNOR2_X1 U652 ( .A(KEYINPUT41), .B(n565), .ZN(n645) );
  INV_X1 U653 ( .A(n645), .ZN(n618) );
  NAND2_X1 U654 ( .A1(n566), .A2(n618), .ZN(n567) );
  XNOR2_X1 U655 ( .A(n567), .B(KEYINPUT42), .ZN(n744) );
  NOR2_X1 U656 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U657 ( .A(n570), .B(KEYINPUT40), .Z(n745) );
  NOR2_X1 U658 ( .A1(n408), .A2(n571), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n572), .A2(n620), .ZN(n573) );
  XNOR2_X1 U660 ( .A(KEYINPUT43), .B(n573), .ZN(n575) );
  NAND2_X1 U661 ( .A1(n575), .A2(n574), .ZN(n694) );
  INV_X1 U662 ( .A(n576), .ZN(n579) );
  NOR2_X1 U663 ( .A1(G898), .A2(n663), .ZN(n725) );
  NAND2_X1 U664 ( .A1(n577), .A2(n725), .ZN(n578) );
  NAND2_X1 U665 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U666 ( .A(KEYINPUT92), .B(n580), .Z(n581) );
  INV_X1 U667 ( .A(KEYINPUT34), .ZN(n584) );
  XNOR2_X1 U668 ( .A(n585), .B(n584), .ZN(n587) );
  NAND2_X1 U669 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U670 ( .A(n588), .B(KEYINPUT35), .ZN(n739) );
  NOR2_X1 U671 ( .A1(n594), .A2(n590), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U673 ( .A1(n639), .A2(n630), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n599), .A2(n596), .ZN(n682) );
  NAND2_X1 U675 ( .A1(n743), .A2(n682), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT44), .ZN(n614) );
  NAND2_X1 U677 ( .A1(n630), .A2(n599), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U679 ( .A(KEYINPUT105), .B(n602), .Z(n741) );
  XOR2_X1 U680 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n607) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n642) );
  NAND2_X1 U682 ( .A1(n642), .A2(n605), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n607), .B(n606), .ZN(n690) );
  NOR2_X1 U684 ( .A1(n639), .A2(n610), .ZN(n675) );
  NOR2_X1 U685 ( .A1(n690), .A2(n675), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n624), .A2(n611), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n741), .A2(n612), .ZN(n613) );
  INV_X1 U688 ( .A(n615), .ZN(n721) );
  AND2_X1 U689 ( .A1(n617), .A2(n618), .ZN(n652) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n626) );
  NOR2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U694 ( .A1(n628), .A2(n627), .ZN(n647) );
  NOR2_X1 U695 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U696 ( .A(KEYINPUT49), .B(n631), .ZN(n637) );
  NAND2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n635) );
  XOR2_X1 U698 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n634) );
  XNOR2_X1 U699 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U700 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U701 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U702 ( .A(n640), .B(KEYINPUT118), .ZN(n641) );
  NOR2_X1 U703 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U704 ( .A(KEYINPUT51), .B(n643), .Z(n644) );
  NOR2_X1 U705 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U706 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U707 ( .A(n648), .B(KEYINPUT52), .ZN(n649) );
  NOR2_X1 U708 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U709 ( .A1(n652), .A2(n651), .ZN(n653) );
  INV_X1 U710 ( .A(n654), .ZN(n656) );
  NAND2_X1 U711 ( .A1(n656), .A2(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U712 ( .A1(n712), .A2(G210), .ZN(n662) );
  XOR2_X1 U713 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n659) );
  XNOR2_X1 U714 ( .A(n662), .B(n661), .ZN(n665) );
  NOR2_X1 U715 ( .A1(G952), .A2(n663), .ZN(n664) );
  NAND2_X1 U716 ( .A1(n665), .A2(n705), .ZN(n667) );
  INV_X1 U717 ( .A(KEYINPUT56), .ZN(n666) );
  XNOR2_X1 U718 ( .A(n667), .B(n666), .ZN(G51) );
  NAND2_X1 U719 ( .A1(n712), .A2(G472), .ZN(n671) );
  XOR2_X1 U720 ( .A(KEYINPUT62), .B(KEYINPUT88), .Z(n668) );
  XNOR2_X1 U721 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U722 ( .A1(n672), .A2(n705), .ZN(n673) );
  XNOR2_X1 U723 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U724 ( .A1(n687), .A2(n675), .ZN(n674) );
  XNOR2_X1 U725 ( .A(G104), .B(n674), .ZN(G6) );
  XOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n677) );
  NAND2_X1 U727 ( .A1(n675), .A2(n689), .ZN(n676) );
  XNOR2_X1 U728 ( .A(n677), .B(n676), .ZN(n678) );
  XOR2_X1 U729 ( .A(n678), .B(KEYINPUT111), .Z(n680) );
  XNOR2_X1 U730 ( .A(G107), .B(KEYINPUT26), .ZN(n679) );
  XNOR2_X1 U731 ( .A(n680), .B(n679), .ZN(G9) );
  XOR2_X1 U732 ( .A(G110), .B(KEYINPUT113), .Z(n681) );
  XNOR2_X1 U733 ( .A(n682), .B(n681), .ZN(G12) );
  XOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .Z(n684) );
  NAND2_X1 U735 ( .A1(n351), .A2(n689), .ZN(n683) );
  XNOR2_X1 U736 ( .A(n684), .B(n683), .ZN(G30) );
  NAND2_X1 U737 ( .A1(n351), .A2(n687), .ZN(n685) );
  XNOR2_X1 U738 ( .A(n685), .B(KEYINPUT114), .ZN(n686) );
  XNOR2_X1 U739 ( .A(G146), .B(n686), .ZN(G48) );
  NAND2_X1 U740 ( .A1(n690), .A2(n687), .ZN(n688) );
  XNOR2_X1 U741 ( .A(n688), .B(G113), .ZN(G15) );
  NAND2_X1 U742 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n691), .B(G116), .ZN(G18) );
  XOR2_X1 U744 ( .A(G134), .B(n692), .Z(n693) );
  XNOR2_X1 U745 ( .A(KEYINPUT116), .B(n693), .ZN(G36) );
  XNOR2_X1 U746 ( .A(G140), .B(n694), .ZN(G42) );
  INV_X1 U747 ( .A(n705), .ZN(n716) );
  XNOR2_X1 U748 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n697) );
  XNOR2_X1 U749 ( .A(n695), .B(KEYINPUT57), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U751 ( .A1(n712), .A2(G469), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n716), .A2(n700), .ZN(G54) );
  NAND2_X1 U754 ( .A1(G475), .A2(n712), .ZN(n704) );
  XNOR2_X1 U755 ( .A(n701), .B(KEYINPUT66), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U758 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(G60) );
  NAND2_X1 U760 ( .A1(G478), .A2(n712), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U762 ( .A1(n716), .A2(n711), .ZN(G63) );
  NAND2_X1 U763 ( .A1(G217), .A2(n712), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U765 ( .A1(n716), .A2(n715), .ZN(G66) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n717), .B(KEYINPUT61), .ZN(n718) );
  XNOR2_X1 U768 ( .A(KEYINPUT122), .B(n718), .ZN(n719) );
  NAND2_X1 U769 ( .A1(n719), .A2(G898), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n720), .B(KEYINPUT123), .ZN(n723) );
  NOR2_X1 U771 ( .A1(n721), .A2(G953), .ZN(n722) );
  NOR2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U773 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U774 ( .A(n727), .B(n726), .Z(G69) );
  XNOR2_X1 U775 ( .A(KEYINPUT124), .B(n728), .ZN(n730) );
  XNOR2_X1 U776 ( .A(n730), .B(n729), .ZN(n732) );
  NOR2_X1 U777 ( .A1(G953), .A2(n731), .ZN(n737) );
  XNOR2_X1 U778 ( .A(n732), .B(KEYINPUT125), .ZN(n733) );
  XNOR2_X1 U779 ( .A(G227), .B(n733), .ZN(n735) );
  NAND2_X1 U780 ( .A1(G900), .A2(G953), .ZN(n734) );
  NOR2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U782 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U783 ( .A(KEYINPUT126), .B(n738), .ZN(G72) );
  XNOR2_X1 U784 ( .A(G122), .B(n739), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n740), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U786 ( .A(G101), .B(n741), .Z(G3) );
  XNOR2_X1 U787 ( .A(G125), .B(n742), .ZN(G27) );
  XNOR2_X1 U788 ( .A(G119), .B(n743), .ZN(G21) );
  XNOR2_X1 U789 ( .A(G137), .B(n744), .ZN(G39) );
  XNOR2_X1 U790 ( .A(G131), .B(n745), .ZN(G33) );
  XNOR2_X1 U791 ( .A(n746), .B(G143), .ZN(G45) );
endmodule

