//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n215), .A2(G50), .A3(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n209), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G107), .ZN(new_n231));
  INV_X1    g0031(.A(G264), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n211), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n214), .B(new_n221), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n235), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G58), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n223), .ZN(new_n256));
  OAI21_X1  g0056(.A(G20), .B1(new_n256), .B2(new_n201), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G159), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT7), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n262), .A2(new_n263), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT7), .B1(new_n269), .B2(new_n209), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(KEYINPUT16), .B(new_n261), .C1(new_n271), .C2(new_n223), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT16), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n263), .B1(new_n262), .B2(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n223), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n273), .B1(new_n276), .B2(new_n260), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n219), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n272), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT68), .ZN(new_n282));
  INV_X1    g0082(.A(new_n279), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G1), .B2(new_n209), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n294), .A3(G274), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(G232), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n266), .A2(new_n268), .A3(G226), .A4(G1698), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G87), .ZN(new_n300));
  OR2_X1    g0100(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n301), .A2(new_n266), .A3(new_n268), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G223), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n299), .B(new_n300), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n294), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(G169), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n289), .A2(KEYINPUT18), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT18), .B1(new_n289), .B2(new_n311), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI211_X1 g0117(.A(KEYINPUT75), .B(KEYINPUT18), .C1(new_n289), .C2(new_n311), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT76), .ZN(new_n321));
  INV_X1    g0121(.A(G200), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n307), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  AOI211_X1 g0124(.A(new_n324), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n307), .A2(G190), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(KEYINPUT76), .C1(new_n322), .C2(new_n307), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n280), .A2(new_n288), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT17), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n320), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT10), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n306), .A2(new_n292), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT66), .B(G226), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n295), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT67), .B(G1698), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n269), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G222), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n262), .A2(G1698), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(new_n229), .B2(new_n262), .C1(new_n304), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n338), .B1(new_n343), .B2(new_n306), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G190), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n282), .A2(new_n209), .A3(G33), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n283), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n283), .A3(new_n286), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G50), .B2(new_n286), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n345), .B1(new_n322), .B2(new_n344), .C1(KEYINPUT9), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n353), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT73), .B(new_n334), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n344), .A2(new_n322), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G190), .B2(new_n344), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n353), .B2(KEYINPUT9), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n356), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n360), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n355), .B1(G169), .B2(new_n344), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n344), .A2(new_n308), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n358), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  INV_X1    g0170(.A(G226), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n370), .B1(new_n303), .B2(new_n371), .C1(new_n240), .C2(new_n342), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n306), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n374));
  INV_X1    g0174(.A(new_n295), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G238), .B2(new_n335), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n373), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g0178(.A(G169), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n373), .A2(new_n376), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT13), .ZN(new_n383));
  OAI211_X1 g0183(.A(G179), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(G169), .C1(new_n377), .C2(new_n378), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n380), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n223), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n209), .A2(G33), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n229), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n279), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT11), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n391), .A2(new_n392), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT12), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n287), .B2(new_n223), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n286), .A2(KEYINPUT12), .A3(G68), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n284), .A2(new_n223), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n394), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n387), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(G190), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n377), .B2(new_n378), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n400), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n342), .A2(new_n224), .B1(new_n231), .B2(new_n262), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT70), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n303), .B2(new_n240), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n340), .A2(KEYINPUT70), .A3(G232), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(new_n294), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n375), .B1(G244), .B2(new_n335), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n308), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n284), .A2(new_n229), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n416), .A2(new_n389), .B1(new_n209), .B2(new_n229), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT71), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n281), .B(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n258), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n415), .B1(G77), .B2(new_n286), .C1(new_n420), .C2(new_n283), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n413), .B1(new_n411), .B2(new_n294), .ZN(new_n422));
  INV_X1    g0222(.A(G169), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n414), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n412), .A2(G190), .A3(new_n413), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n421), .B1(G200), .B2(new_n422), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT72), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n422), .A2(G200), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n420), .A2(new_n283), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n415), .B1(G77), .B2(new_n286), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(KEYINPUT72), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n425), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NOR4_X1   g0236(.A1(new_n333), .A2(new_n369), .A3(new_n406), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT81), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT80), .ZN(new_n440));
  AND2_X1   g0240(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n262), .A3(G244), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT4), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(KEYINPUT77), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n266), .A2(new_n268), .A3(G250), .A4(G1698), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n262), .A2(KEYINPUT79), .A3(G250), .A4(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT77), .B1(new_n444), .B2(new_n445), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n443), .A2(new_n262), .A3(KEYINPUT4), .A4(G244), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n294), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n208), .A2(G45), .ZN(new_n463));
  OR2_X1    g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n306), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G257), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n294), .A2(G274), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n440), .B1(new_n462), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n454), .A2(new_n459), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n445), .B1(new_n303), .B2(new_n230), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n474), .A2(new_n477), .A3(new_n446), .A4(new_n451), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n306), .ZN(new_n479));
  INV_X1    g0279(.A(new_n472), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(KEYINPUT80), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(G169), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n231), .A2(KEYINPUT6), .A3(G97), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n231), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n205), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(KEYINPUT6), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n271), .B2(new_n231), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n279), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n287), .A2(new_n484), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n208), .A2(G33), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n283), .A2(new_n286), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(new_n484), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n479), .A2(new_n480), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G179), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n439), .B1(new_n482), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT80), .B1(new_n479), .B2(new_n480), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n440), .B(new_n472), .C1(new_n478), .C2(new_n306), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n423), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n462), .A2(new_n472), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(new_n308), .B1(new_n490), .B2(new_n495), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n496), .B1(G200), .B2(new_n497), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n473), .A2(new_n481), .A3(G190), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n499), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT86), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n466), .A2(new_n306), .A3(new_n232), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n262), .A2(G257), .A3(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n513), .C1(new_n226), .C2(new_n303), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(new_n306), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n308), .A3(new_n471), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n306), .ZN(new_n517));
  INV_X1    g0317(.A(new_n511), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n517), .A2(new_n471), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n516), .B1(new_n519), .B2(G169), .ZN(new_n520));
  INV_X1    g0320(.A(new_n493), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT25), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n286), .B2(G107), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n287), .A2(KEYINPUT25), .A3(new_n231), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n521), .A2(G107), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n266), .A2(new_n268), .A3(new_n209), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n262), .A2(new_n529), .A3(new_n209), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(G20), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n209), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n231), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n531), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n526), .B1(new_n542), .B2(new_n279), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n510), .B1(new_n520), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n515), .A2(new_n471), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n543), .B(new_n546), .C1(new_n324), .C2(new_n545), .ZN(new_n547));
  INV_X1    g0347(.A(new_n541), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n540), .B1(new_n531), .B2(new_n537), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n279), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n525), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n545), .A2(new_n423), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(KEYINPUT86), .A3(new_n552), .A4(new_n516), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n544), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n467), .A2(G270), .B1(new_n470), .B2(new_n466), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n266), .A2(new_n268), .A3(G257), .ZN(new_n556));
  INV_X1    g0356(.A(G303), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n556), .A2(new_n339), .B1(new_n262), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n262), .A2(G264), .A3(G1698), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n306), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n423), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  INV_X1    g0363(.A(G116), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n287), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n493), .B2(new_n564), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT20), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n209), .B1(new_n484), .B2(G33), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n457), .B2(new_n458), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n278), .A2(new_n219), .B1(G20), .B2(new_n564), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n458), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n456), .ZN(new_n574));
  OAI211_X1 g0374(.A(KEYINPUT20), .B(new_n570), .C1(new_n574), .C2(new_n568), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n566), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n562), .A2(new_n563), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n576), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT21), .B1(new_n578), .B2(new_n561), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n209), .B1(new_n370), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G87), .B2(new_n206), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n266), .A2(new_n268), .A3(new_n209), .A4(G68), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n585), .A2(KEYINPUT82), .A3(new_n581), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT82), .B1(new_n585), .B2(new_n581), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n583), .B(new_n584), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n279), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n416), .A2(new_n287), .ZN(new_n590));
  INV_X1    g0390(.A(new_n416), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n521), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT83), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n588), .A2(new_n279), .B1(new_n287), .B2(new_n416), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n294), .A2(G250), .A3(new_n463), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n469), .B2(new_n463), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(G1698), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n532), .B(new_n601), .C1(new_n303), .C2(new_n224), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n600), .B1(new_n602), .B2(new_n306), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(G169), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n308), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(G190), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n521), .A2(G87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n589), .A2(new_n590), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n602), .A2(new_n306), .ZN(new_n609));
  INV_X1    g0409(.A(new_n600), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n322), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n598), .A2(new_n605), .B1(new_n606), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n555), .A2(new_n560), .A3(G179), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n576), .A3(KEYINPUT84), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT84), .B1(new_n614), .B2(new_n576), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT85), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n555), .A2(new_n560), .A3(G190), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n576), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n322), .B1(new_n555), .B2(new_n560), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n622), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT85), .A3(new_n576), .A4(new_n620), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n580), .A2(new_n613), .A3(new_n618), .A4(new_n626), .ZN(new_n627));
  NOR4_X1   g0427(.A1(new_n438), .A2(new_n509), .A3(new_n554), .A4(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n368), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n316), .A2(new_n312), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n332), .A2(new_n405), .ZN(new_n631));
  INV_X1    g0431(.A(new_n425), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n387), .B2(new_n401), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n358), .A2(new_n365), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n482), .A2(new_n498), .ZN(new_n637));
  INV_X1    g0437(.A(new_n606), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n595), .B(new_n607), .C1(new_n603), .C2(new_n322), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n598), .B2(new_n605), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT26), .B1(new_n637), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n613), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n499), .B2(new_n505), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n644), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n598), .A2(new_n605), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n563), .B1(new_n562), .B2(new_n576), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n578), .A2(KEYINPUT21), .A3(new_n561), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  INV_X1    g0451(.A(new_n614), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n578), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n649), .B(new_n650), .C1(new_n653), .C2(new_n615), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n520), .A2(new_n543), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n643), .B(new_n547), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n648), .B1(new_n509), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n636), .B1(new_n438), .B2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  INV_X1    g0460(.A(new_n626), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n654), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT88), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT27), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT88), .A4(G13), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G213), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n663), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n671), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(KEYINPUT89), .A3(G213), .A4(new_n669), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n578), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n580), .A2(new_n618), .A3(new_n626), .A4(KEYINPUT90), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n662), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n654), .A2(new_n678), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G330), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n677), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n543), .ZN(new_n685));
  INV_X1    g0485(.A(new_n655), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n554), .A2(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n654), .A2(new_n684), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n677), .B(new_n690), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n554), .A2(new_n689), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n212), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n217), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  INV_X1    g0501(.A(new_n648), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n643), .A2(new_n502), .A3(new_n504), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(KEYINPUT26), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n544), .A2(new_n553), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n547), .B(new_n643), .C1(new_n705), .C2(new_n654), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n509), .B2(new_n706), .ZN(new_n707));
  AOI211_X1 g0507(.A(KEYINPUT26), .B(new_n645), .C1(new_n499), .C2(new_n505), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT29), .B(new_n684), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n499), .A2(new_n505), .A3(new_n508), .ZN(new_n710));
  INV_X1    g0510(.A(new_n656), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n702), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n482), .A2(new_n498), .A3(new_n439), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT81), .B1(new_n502), .B2(new_n504), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT26), .B(new_n613), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n644), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n691), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n709), .B1(new_n718), .B2(KEYINPUT29), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n652), .A2(new_n515), .A3(new_n603), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(new_n473), .A3(new_n481), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n720), .A2(new_n473), .A3(new_n481), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n603), .A2(G179), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n555), .A2(new_n560), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n545), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n503), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n722), .B2(new_n724), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n684), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n627), .A2(new_n554), .ZN(new_n737));
  INV_X1    g0537(.A(new_n691), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n710), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n719), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n701), .B1(new_n743), .B2(G1), .ZN(G364));
  AND2_X1   g0544(.A1(new_n209), .A2(G13), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n208), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n696), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n683), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n680), .A2(new_n681), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT99), .Z(new_n756));
  OR2_X1    g0556(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n212), .A2(new_n262), .ZN(new_n758));
  INV_X1    g0558(.A(G355), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(G116), .B2(new_n212), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n695), .A2(new_n262), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n218), .B2(new_n291), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n250), .A2(new_n291), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n219), .B1(G20), .B2(new_n423), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n748), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT95), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n209), .A2(new_n308), .A3(new_n322), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n770), .B1(new_n774), .B2(G190), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n772), .A2(KEYINPUT95), .A3(new_n324), .A4(new_n773), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n209), .A2(new_n324), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n308), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n777), .A2(new_n778), .B1(G322), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n774), .A2(new_n324), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G326), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n209), .B1(new_n787), .B2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(G294), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n209), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n780), .A2(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n269), .B1(new_n788), .B2(new_n789), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n322), .A2(G179), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT96), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n791), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n791), .A2(new_n787), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G283), .A2(new_n799), .B1(new_n801), .B2(G329), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n797), .A2(new_n557), .B1(KEYINPUT97), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n793), .B(new_n804), .C1(KEYINPUT97), .C2(new_n803), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n784), .A2(new_n786), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n777), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n223), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n262), .B1(new_n795), .B2(new_n225), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT94), .Z(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G50), .B2(new_n785), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n781), .A2(new_n255), .B1(new_n792), .B2(new_n229), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT92), .Z(new_n813));
  NOR2_X1   g0613(.A1(new_n788), .A2(new_n484), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G107), .B2(new_n799), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n801), .A2(G159), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT32), .Z(new_n817));
  NAND4_X1  g0617(.A1(new_n811), .A2(new_n813), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n806), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n769), .B1(new_n819), .B2(new_n766), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n749), .A2(new_n752), .B1(new_n757), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NOR2_X1   g0622(.A1(new_n425), .A2(new_n677), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n684), .A2(new_n433), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n429), .B2(new_n435), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n691), .B(new_n823), .C1(new_n826), .C2(new_n425), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n647), .B2(new_n657), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n823), .B1(new_n826), .B2(new_n425), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n718), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n748), .B1(new_n830), .B2(new_n741), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n741), .B2(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(new_n785), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n833), .A2(new_n557), .B1(new_n564), .B2(new_n792), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n777), .B2(G283), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT102), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n797), .A2(new_n231), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G294), .A2(new_n782), .B1(new_n801), .B2(G311), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(new_n269), .C1(new_n225), .C2(new_n798), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n836), .A2(new_n814), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n792), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G143), .A2(new_n782), .B1(new_n841), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n833), .C1(new_n807), .C2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n797), .A2(new_n202), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n269), .B1(new_n799), .B2(G68), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n255), .B2(new_n788), .C1(new_n851), .C2(new_n800), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n766), .B1(new_n840), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n766), .A2(new_n753), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT100), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n748), .B1(new_n856), .B2(G77), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT101), .Z(new_n858));
  OAI211_X1 g0658(.A(new_n854), .B(new_n858), .C1(new_n829), .C2(new_n754), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n832), .A2(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n745), .A2(new_n208), .ZN(new_n861));
  INV_X1    g0661(.A(G330), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n330), .A2(new_n675), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n315), .B1(new_n313), .B2(new_n312), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n318), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n289), .B1(new_n326), .B2(new_n328), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT17), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT17), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n331), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n289), .A2(new_n311), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n331), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n863), .B1(new_n874), .B2(KEYINPUT105), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT105), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n331), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n872), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n672), .A2(new_n674), .A3(KEYINPUT107), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT107), .B1(new_n672), .B2(new_n674), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT37), .B1(new_n883), .B2(new_n289), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n289), .A2(KEYINPUT106), .A3(new_n311), .ZN(new_n885));
  AND4_X1   g0685(.A1(new_n331), .A2(new_n880), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n871), .B(KEYINPUT38), .C1(new_n878), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n289), .A2(new_n311), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT108), .B1(new_n866), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n883), .A2(new_n289), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT108), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n331), .A2(new_n892), .A3(new_n873), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n886), .B1(new_n894), .B2(KEYINPUT37), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n891), .B1(new_n332), .B2(new_n630), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n739), .A2(new_n735), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n823), .ZN(new_n901));
  INV_X1    g0701(.A(new_n426), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(KEYINPUT72), .B2(new_n434), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n427), .A2(new_n428), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n824), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n905), .B2(new_n632), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n401), .A2(new_n677), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n402), .A2(new_n405), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n405), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n401), .B(new_n677), .C1(new_n387), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n906), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n898), .A2(new_n900), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n900), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT105), .B1(new_n866), .B2(new_n889), .ZN(new_n915));
  INV_X1    g0715(.A(new_n863), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n877), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n886), .B1(new_n917), .B2(KEYINPUT37), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n320), .B2(new_n332), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n888), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n887), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n912), .A2(KEYINPUT40), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT109), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n739), .A2(new_n735), .A3(new_n899), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n438), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n862), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n923), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n630), .A2(new_n883), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n920), .A2(new_n887), .A3(KEYINPUT39), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT39), .B1(new_n887), .B2(new_n897), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n387), .A2(new_n401), .A3(new_n684), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n928), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n908), .A2(new_n910), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n826), .A2(new_n425), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n738), .A3(new_n901), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n712), .B2(new_n717), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT104), .B1(new_n939), .B2(new_n823), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT104), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n828), .A2(new_n941), .A3(new_n901), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n936), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n921), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n636), .B1(new_n719), .B2(new_n438), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n861), .B1(new_n927), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n927), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n220), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT36), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n217), .A2(new_n229), .A3(new_n256), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n202), .B2(G68), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n955), .A2(new_n208), .A3(G13), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT103), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n953), .A3(new_n957), .ZN(G367));
  OR2_X1    g0758(.A1(new_n554), .A2(new_n689), .ZN(new_n959));
  INV_X1    g0759(.A(new_n689), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n687), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT110), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n682), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n682), .A2(new_n962), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n680), .A2(KEYINPUT110), .A3(G330), .A4(new_n681), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n719), .A3(new_n741), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT111), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n691), .A2(new_n496), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n499), .A2(new_n505), .A3(new_n508), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n637), .A2(new_n691), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n693), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n693), .A3(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n974), .B2(new_n693), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n692), .A2(new_n972), .A3(KEYINPUT44), .A4(new_n973), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n979), .A2(new_n688), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n688), .B1(new_n979), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n967), .A2(new_n719), .A3(new_n741), .A4(KEYINPUT111), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n970), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT112), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT112), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n970), .A2(new_n986), .A3(new_n990), .A4(new_n987), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n742), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n696), .B(KEYINPUT41), .Z(new_n993));
  OAI21_X1  g0793(.A(new_n746), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n959), .B1(new_n972), .B2(new_n973), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n974), .A2(new_n705), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n499), .A2(new_n505), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n738), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n677), .A2(new_n608), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n643), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n648), .B2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n996), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n683), .A2(new_n687), .A3(new_n974), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n796), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n798), .A2(new_n484), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G317), .B2(new_n801), .ZN(new_n1011));
  INV_X1    g0811(.A(G283), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n792), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n795), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(G116), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n269), .B1(new_n788), .B2(new_n231), .C1(new_n557), .C2(new_n781), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1009), .A2(new_n1013), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n789), .B2(new_n807), .C1(new_n790), .C2(new_n833), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n262), .B1(new_n798), .B2(new_n229), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n788), .A2(new_n223), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n781), .A2(new_n844), .B1(new_n792), .B2(new_n202), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n795), .A2(new_n255), .B1(new_n800), .B2(new_n843), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n785), .A2(G143), .ZN(new_n1026));
  INV_X1    g0826(.A(G159), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1026), .C1(new_n1027), .C2(new_n807), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1019), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT47), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n766), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n768), .B1(new_n695), .B2(new_n591), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n761), .A2(new_n246), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n696), .B(new_n747), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1031), .B(new_n1034), .C1(new_n756), .C2(new_n1002), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1008), .A2(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n970), .A2(new_n987), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n696), .C1(new_n743), .C2(new_n967), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n967), .A2(new_n747), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n758), .A2(new_n698), .B1(G107), .B2(new_n212), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n698), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT115), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n291), .B1(new_n223), .B2(new_n229), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT116), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n419), .A2(new_n202), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT117), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT50), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n762), .B1(new_n243), .B2(G45), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1040), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n748), .B1(new_n1052), .B2(new_n768), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G50), .A2(new_n782), .B1(new_n801), .B2(G150), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n223), .B2(new_n792), .C1(new_n229), .C2(new_n795), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n788), .A2(new_n416), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1055), .A2(new_n269), .A3(new_n1010), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n777), .A2(new_n282), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n785), .A2(KEYINPUT118), .A3(G159), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT118), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n833), .B2(new_n1027), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n262), .B1(new_n801), .B2(G326), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n795), .A2(new_n789), .B1(new_n788), .B2(new_n1012), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G317), .A2(new_n782), .B1(new_n841), .B2(G303), .ZN(new_n1065));
  INV_X1    g0865(.A(G322), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n833), .C1(new_n807), .C2(new_n790), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1063), .B1(new_n564), .B2(new_n798), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1062), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1053), .B1(new_n1074), .B2(new_n766), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n687), .B2(new_n756), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1038), .A2(new_n1039), .A3(new_n1076), .ZN(G393));
  NAND3_X1  g0877(.A1(new_n972), .A2(new_n755), .A3(new_n973), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n788), .A2(new_n229), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G68), .A2(new_n1015), .B1(new_n801), .B2(G143), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n262), .C1(new_n225), .C2(new_n798), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(new_n419), .C2(new_n841), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n202), .B2(new_n807), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n785), .A2(G150), .B1(G159), .B2(new_n782), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n785), .A2(G317), .B1(G311), .B2(new_n782), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n795), .A2(new_n1012), .B1(new_n800), .B2(new_n1066), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n269), .B1(new_n788), .B2(new_n564), .C1(new_n231), .C2(new_n798), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G294), .C2(new_n841), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n807), .B2(new_n557), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1083), .A2(new_n1085), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n766), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n767), .B1(new_n484), .B2(new_n212), .C1(new_n762), .C2(new_n253), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1078), .A2(new_n748), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n986), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n746), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n989), .A2(new_n991), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n697), .B1(new_n1037), .B2(new_n1096), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  NAND2_X1  g0901(.A1(new_n935), .A2(new_n829), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n924), .A2(new_n862), .A3(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n828), .A2(new_n941), .A3(new_n901), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n941), .B1(new_n828), .B2(new_n901), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n935), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n931), .B1(new_n1106), .B2(new_n932), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n684), .B(new_n937), .C1(new_n707), .C2(new_n708), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n901), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n932), .B(new_n898), .C1(new_n1110), .C2(new_n936), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1103), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n943), .A2(new_n933), .B1(new_n930), .B2(new_n929), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n862), .B1(new_n736), .B2(new_n739), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n829), .A3(new_n935), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n924), .A2(new_n862), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n437), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n636), .C1(new_n438), .C2(new_n719), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n935), .B1(new_n1115), .B2(new_n829), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1122), .A2(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n900), .A2(G330), .A3(new_n829), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n936), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1116), .A2(new_n1125), .A3(new_n1110), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1121), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1113), .A2(new_n1117), .A3(new_n1127), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n696), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1113), .A2(new_n1117), .A3(new_n747), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n748), .B1(new_n856), .B2(new_n282), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n781), .A2(new_n564), .B1(new_n792), .B2(new_n484), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n269), .B1(new_n788), .B2(new_n229), .C1(new_n223), .C2(new_n798), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(G294), .C2(new_n801), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n225), .B2(new_n797), .C1(new_n1012), .C2(new_n833), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n807), .A2(new_n231), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n785), .A2(G128), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n792), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n798), .A2(new_n202), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G125), .C2(new_n801), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n262), .B1(new_n781), .B2(new_n851), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n788), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(G159), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n795), .A2(new_n844), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1139), .A2(new_n1143), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n807), .A2(new_n843), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1137), .A2(new_n1138), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1133), .B1(new_n1151), .B2(new_n766), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT119), .Z(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n931), .B2(new_n754), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1132), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1131), .A2(new_n1156), .ZN(G378));
  OAI21_X1  g0957(.A(new_n748), .B1(new_n856), .B2(G50), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n262), .A2(G41), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G50), .B(new_n1159), .C1(new_n265), .C2(new_n290), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n229), .B2(new_n795), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n416), .A2(new_n792), .B1(new_n798), .B2(new_n255), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n781), .A2(new_n231), .B1(new_n800), .B2(new_n1012), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1022), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n564), .B2(new_n833), .C1(new_n807), .C2(new_n484), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT58), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n788), .A2(new_n844), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n782), .A2(G128), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n843), .B2(new_n792), .C1(new_n795), .C2(new_n1140), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(G125), .C2(new_n785), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n851), .B2(new_n807), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n265), .B(new_n290), .C1(new_n798), .C2(new_n1027), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G124), .B2(new_n801), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1158), .B1(new_n1178), .B2(new_n766), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n353), .A2(new_n675), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n369), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n369), .A2(new_n1180), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1179), .B1(new_n1187), .B2(new_n754), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT120), .Z(new_n1189));
  AND2_X1   g0989(.A1(new_n887), .A2(new_n897), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n900), .A2(new_n911), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT40), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n899), .A2(new_n735), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1102), .B1(new_n1193), .B2(new_n739), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n913), .A3(new_n921), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1187), .B1(new_n1196), .B2(G330), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n862), .B(new_n1186), .C1(new_n1192), .C2(new_n1195), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n945), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1186), .B1(new_n922), .B2(new_n862), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1194), .A2(new_n913), .A3(new_n921), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n913), .B1(new_n1194), .B2(new_n898), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1187), .B(G330), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n944), .A3(new_n934), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1189), .B1(new_n1205), .B2(new_n747), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1121), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1130), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n696), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1208), .B2(new_n1205), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1212), .B2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n936), .A2(new_n753), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n748), .B1(new_n856), .B2(G68), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n781), .A2(new_n1012), .B1(new_n792), .B2(new_n231), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n269), .B1(new_n788), .B2(new_n416), .C1(new_n229), .C2(new_n798), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G303), .C2(new_n801), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n484), .B2(new_n797), .C1(new_n789), .C2(new_n833), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n807), .A2(new_n564), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n781), .A2(new_n843), .B1(new_n792), .B2(new_n844), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n262), .B1(new_n788), .B2(new_n202), .C1(new_n255), .C2(new_n798), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G128), .C2(new_n801), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n1027), .B2(new_n797), .C1(new_n851), .C2(new_n833), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n807), .A2(new_n1140), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1221), .A2(new_n1222), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1217), .B1(new_n1228), .B2(new_n766), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1215), .A2(new_n747), .B1(new_n1216), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n993), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1128), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1215), .A2(new_n1207), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  NOR4_X1   g1034(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n697), .B1(new_n1118), .B2(new_n1128), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1155), .B1(new_n1236), .B2(new_n1130), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1235), .A2(new_n1100), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G375), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1238), .A2(new_n1008), .A3(new_n1035), .A4(new_n1239), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n676), .A2(G213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1237), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1206), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1208), .A2(new_n1231), .A3(new_n1205), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1205), .A2(new_n747), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1188), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1237), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1242), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1123), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n1126), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(new_n696), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1127), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1255), .B2(new_n1233), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(G384), .A3(new_n1230), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1256), .B2(new_n1230), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1251), .A2(KEYINPUT62), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1260), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1251), .A2(new_n1260), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1267));
  XOR2_X1   g1067(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1268));
  NAND2_X1  g1068(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1241), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1242), .A2(G2897), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT121), .Z(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1259), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1257), .A3(new_n1272), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1268), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1267), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1245), .B1(new_n1264), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(new_n1100), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(new_n821), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1008), .A2(new_n1035), .A3(G390), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1282), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G390), .B1(new_n1008), .B2(new_n1035), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1035), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1287), .B(new_n1100), .C1(new_n994), .C2(new_n1007), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1285), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1251), .A2(KEYINPUT62), .A3(new_n1260), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(KEYINPUT126), .A3(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1267), .A4(new_n1278), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1280), .A2(new_n1290), .A3(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1241), .A4(new_n1260), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT123), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1251), .A2(KEYINPUT123), .A3(KEYINPUT63), .A4(new_n1260), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1270), .A2(KEYINPUT122), .A3(new_n1277), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT122), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1251), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT63), .B1(new_n1251), .B2(new_n1260), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1284), .A2(new_n1289), .A3(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(new_n1305), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT124), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1300), .A2(new_n1305), .A3(new_n1309), .A4(KEYINPUT124), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1295), .A2(new_n1314), .ZN(G405));
  NOR2_X1   g1115(.A1(new_n1239), .A2(G378), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1246), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  XOR2_X1   g1118(.A(new_n1318), .B(new_n1260), .Z(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1290), .ZN(G402));
endmodule


