//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1143, new_n1144, new_n1145, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT68), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND4_X1  g037(.A1(new_n459), .A2(new_n461), .A3(G137), .A4(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n458), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT72), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n460), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT69), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g056(.A(KEYINPUT71), .B(G2105), .C1(new_n475), .C2(new_n478), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n468), .B1(new_n481), .B2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n459), .A2(new_n461), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT73), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT73), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n459), .A2(new_n461), .A3(new_n486), .A4(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n484), .A2(KEYINPUT74), .A3(new_n462), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT74), .B1(new_n484), .B2(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NOR2_X1   g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n489), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  NOR2_X1   g072(.A1(KEYINPUT4), .A2(G2105), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT69), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT69), .B1(new_n459), .B2(new_n461), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n459), .A2(new_n461), .A3(G138), .A4(new_n462), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G114), .A2(G2104), .ZN(new_n508));
  INV_X1    g083(.A(G126), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n484), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G2105), .B1(G102), .B2(new_n465), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n507), .A2(KEYINPUT76), .A3(new_n511), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n525), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  AOI22_X1  g108(.A1(new_n526), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n534));
  INV_X1    g109(.A(new_n522), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n529), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n536), .B1(G51), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n537), .A2(G52), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OAI221_X1 g120(.A(new_n543), .B1(new_n544), .B2(new_n527), .C1(new_n545), .C2(new_n524), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(new_n527), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G81), .B1(G43), .B2(new_n537), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n524), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n537), .A2(KEYINPUT77), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n561), .A4(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n535), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n560), .A2(new_n562), .B1(G651), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n548), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(new_n537), .A2(G49), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT78), .Z(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n548), .A2(G87), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n548), .A2(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n537), .A2(G48), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT79), .Z(new_n577));
  AND3_X1   g152(.A1(new_n519), .A2(new_n521), .A3(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n524), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT80), .B(G47), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n527), .A2(new_n583), .B1(new_n529), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n522), .A2(G92), .A3(new_n526), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  AOI22_X1  g165(.A1(new_n522), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n524), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n537), .A2(G54), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n588), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n588), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n606), .B(new_n607), .C1(G868), .C2(new_n552), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g184(.A1(new_n499), .A2(new_n500), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n465), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n492), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n488), .A2(G135), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n619), .B(new_n620), .C1(G111), .C2(new_n462), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT83), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2443), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT85), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2430), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2435), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2438), .Z(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n633), .B(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(G14), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT17), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n644), .B2(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2096), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n658), .A2(KEYINPUT87), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(KEYINPUT87), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n655), .A2(new_n656), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n658), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n662), .A2(new_n666), .ZN(new_n669));
  NAND4_X1  g244(.A1(new_n665), .A2(new_n667), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G4), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n595), .B2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(G1348), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(G19), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n552), .B2(new_n677), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1341), .ZN(new_n684));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G26), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n492), .A2(G128), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n488), .A2(G140), .ZN(new_n688));
  OR2_X1    g263(.A1(G104), .A2(G2105), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n689), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n686), .B1(new_n692), .B2(new_n685), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n686), .B(new_n693), .S(KEYINPUT28), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT92), .B(G2067), .Z(new_n695));
  AOI21_X1  g270(.A(new_n684), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n681), .B(new_n696), .C1(new_n695), .C2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n685), .A2(G33), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n611), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(new_n462), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n465), .A2(G103), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT25), .Z(new_n703));
  AND3_X1   g278(.A1(new_n488), .A2(KEYINPUT94), .A3(G139), .ZN(new_n704));
  AOI21_X1  g279(.A(KEYINPUT94), .B1(new_n488), .B2(G139), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n701), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n699), .B1(new_n707), .B2(new_n685), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G2072), .Z(new_n709));
  AOI22_X1  g284(.A1(new_n492), .A2(G129), .B1(G141), .B2(new_n488), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT95), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n465), .A2(G105), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G29), .B2(G32), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  OR2_X1    g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT24), .A2(G34), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n685), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G160), .B2(new_n685), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n718), .A2(new_n719), .B1(new_n723), .B2(G2084), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT96), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n677), .A2(G20), .ZN(new_n727));
  OAI211_X1 g302(.A(KEYINPUT23), .B(new_n727), .C1(new_n599), .C2(new_n677), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(KEYINPUT23), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1956), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n623), .A2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n718), .B2(new_n719), .ZN(new_n732));
  NAND2_X1  g307(.A1(G171), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G5), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT30), .B(G28), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n734), .A2(new_n735), .B1(new_n685), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n735), .B2(new_n734), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G21), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G168), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT97), .B(G1966), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n732), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n723), .A2(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT98), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n730), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n685), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n685), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2090), .ZN(new_n751));
  NOR2_X1   g326(.A1(G27), .A2(G29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G164), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2078), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n726), .A2(new_n747), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n677), .A2(G22), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G166), .B2(new_n677), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1971), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n677), .A2(G23), .ZN(new_n759));
  INV_X1    g334(.A(G288), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n677), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT33), .Z(new_n762));
  AOI21_X1  g337(.A(new_n758), .B1(new_n762), .B2(G1976), .ZN(new_n763));
  MUX2_X1   g338(.A(G6), .B(G305), .S(G16), .Z(new_n764));
  XOR2_X1   g339(.A(KEYINPUT32), .B(G1981), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n766), .C1(G1976), .C2(new_n762), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n685), .A2(G25), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n492), .A2(G119), .ZN(new_n772));
  OAI21_X1  g347(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n773));
  INV_X1    g348(.A(G95), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n462), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n488), .B2(G131), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(new_n685), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT35), .B(G1991), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n677), .A2(G24), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n586), .B2(new_n677), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT88), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1986), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n769), .A2(new_n770), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT91), .Z(new_n789));
  AND3_X1   g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n698), .B(new_n755), .C1(new_n790), .C2(new_n791), .ZN(G150));
  INV_X1    g367(.A(G150), .ZN(G311));
  XOR2_X1   g368(.A(KEYINPUT100), .B(G93), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT99), .B(G55), .Z(new_n795));
  OAI22_X1  g370(.A1(new_n527), .A2(new_n794), .B1(new_n529), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT101), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(new_n524), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G860), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT37), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n552), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT38), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n593), .A2(new_n594), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n602), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n808));
  AOI21_X1  g383(.A(G860), .B1(new_n808), .B2(KEYINPUT102), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(KEYINPUT102), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n810), .B2(new_n811), .ZN(G145));
  XNOR2_X1  g387(.A(G162), .B(G160), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(new_n623), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n692), .A2(new_n715), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n692), .A2(new_n715), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n507), .A2(new_n511), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n817), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n512), .B1(new_n820), .B2(new_n815), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n819), .B2(new_n821), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n707), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n819), .A2(new_n821), .A3(new_n706), .ZN(new_n828));
  OAI211_X1 g403(.A(KEYINPUT104), .B(new_n707), .C1(new_n823), .C2(new_n824), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n492), .A2(G130), .ZN(new_n831));
  OR2_X1    g406(.A1(G106), .A2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n488), .B2(G142), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n613), .B(new_n777), .ZN(new_n838));
  INV_X1    g413(.A(new_n836), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n827), .A2(new_n839), .A3(new_n828), .A4(new_n829), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n838), .B1(new_n837), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n814), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(new_n814), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT40), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n844), .A2(new_n847), .A3(new_n851), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G395));
  XOR2_X1   g428(.A(new_n803), .B(KEYINPUT105), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n604), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n595), .A2(new_n599), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n805), .A2(G299), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT106), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n856), .A2(KEYINPUT41), .A3(new_n857), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(new_n856), .B2(new_n857), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n864), .B1(new_n855), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n870));
  XNOR2_X1  g445(.A(G288), .B(G166), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n586), .ZN(new_n872));
  XNOR2_X1  g447(.A(G288), .B(G303), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G290), .ZN(new_n874));
  XOR2_X1   g449(.A(G305), .B(KEYINPUT107), .Z(new_n875));
  AND3_X1   g450(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n864), .B(new_n879), .C1(new_n855), .C2(new_n868), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n870), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n870), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(G868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n800), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(G868), .B2(new_n884), .ZN(G295));
  OAI21_X1  g460(.A(new_n883), .B1(G868), .B2(new_n884), .ZN(G331));
  INV_X1    g461(.A(new_n878), .ZN(new_n887));
  XNOR2_X1  g462(.A(G171), .B(G286), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n803), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n803), .A2(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(KEYINPUT109), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n803), .A2(new_n892), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(new_n868), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(KEYINPUT108), .A3(new_n890), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n803), .A2(new_n897), .A3(new_n888), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n896), .A2(new_n898), .B1(new_n860), .B2(new_n862), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n887), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n867), .A2(new_n896), .A3(new_n898), .ZN(new_n901));
  INV_X1    g476(.A(new_n894), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n878), .B(new_n901), .C1(new_n902), .C2(new_n858), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n903), .A3(new_n848), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n902), .B2(new_n858), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n887), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n848), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n904), .A2(KEYINPUT110), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n900), .A2(new_n903), .A3(new_n914), .A4(new_n848), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(KEYINPUT43), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT111), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n913), .A2(new_n918), .A3(KEYINPUT43), .A4(new_n915), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(KEYINPUT44), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n912), .B1(new_n920), .B2(new_n921), .ZN(G397));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n512), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n467), .B(KEYINPUT72), .Z(new_n927));
  OAI21_X1  g502(.A(G125), .B1(new_n499), .B2(new_n500), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n462), .B1(new_n928), .B2(new_n477), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(KEYINPUT71), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n480), .B(new_n462), .C1(new_n928), .C2(new_n477), .ZN(new_n931));
  OAI211_X1 g506(.A(G40), .B(new_n927), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n691), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n716), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n715), .A2(G1996), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n778), .A2(new_n780), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n692), .A2(new_n935), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n934), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n934), .B1(new_n716), .B2(new_n936), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n933), .A2(KEYINPUT46), .A3(new_n937), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT46), .B1(new_n933), .B2(new_n937), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n777), .B(new_n780), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT112), .Z(new_n951));
  OAI21_X1  g526(.A(new_n933), .B1(new_n951), .B2(new_n940), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n934), .A2(G1986), .A3(G290), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT48), .Z(new_n954));
  AOI211_X1 g529(.A(new_n944), .B(new_n949), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n932), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n514), .A2(new_n923), .A3(new_n515), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n956), .B(new_n957), .C1(new_n958), .C2(KEYINPUT50), .ZN(new_n959));
  INV_X1    g534(.A(G1956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT57), .B1(G299), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT57), .ZN(new_n964));
  AOI211_X1 g539(.A(KEYINPUT117), .B(new_n964), .C1(new_n566), .C2(new_n567), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n958), .A2(new_n925), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n925), .B(G1384), .C1(new_n507), .C2(new_n511), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n932), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT56), .B(G2072), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n961), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT118), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n512), .A2(new_n975), .A3(new_n923), .ZN(new_n976));
  AND3_X1   g551(.A1(G160), .A2(new_n976), .A3(G40), .ZN(new_n977));
  AOI21_X1  g552(.A(G1348), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n924), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(G40), .A3(G160), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G2067), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n973), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n956), .A2(new_n935), .A3(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(G160), .A2(new_n976), .A3(G40), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(KEYINPUT50), .B2(new_n958), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT118), .B(new_n983), .C1(new_n985), .C2(G1348), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n986), .A3(new_n595), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(KEYINPUT119), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n982), .A2(new_n986), .A3(new_n989), .A4(new_n595), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n961), .A2(new_n971), .ZN(new_n991));
  INV_X1    g566(.A(new_n966), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n972), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n974), .A2(new_n977), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n680), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT118), .B1(new_n997), .B2(new_n983), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n978), .A2(new_n973), .A3(new_n981), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT60), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT60), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n982), .A2(new_n986), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n595), .A3(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT60), .B(new_n805), .C1(new_n998), .C2(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT61), .B1(new_n992), .B2(KEYINPUT122), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n961), .A2(new_n966), .A3(new_n971), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n966), .B1(new_n961), .B2(new_n971), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n993), .A2(new_n972), .A3(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT120), .B(G1996), .Z(new_n1012));
  NAND3_X1  g587(.A1(new_n967), .A2(new_n969), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT58), .B(G1341), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n980), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n967), .A2(new_n969), .A3(KEYINPUT121), .A4(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n552), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1019), .B2(new_n552), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1009), .B(new_n1011), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n995), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2084), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n985), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G40), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n924), .B2(new_n925), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(G160), .C1(new_n958), .C2(new_n925), .ZN(new_n1029));
  INV_X1    g604(.A(new_n741), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G168), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1026), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1041), .A3(G286), .ZN(new_n1042));
  NOR2_X1   g617(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1037), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT124), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n1035), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n967), .A2(new_n969), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(G2078), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n996), .A2(new_n735), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n968), .A2(new_n468), .A3(new_n929), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1054), .A2(G2078), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n1028), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n516), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1063), .A2(G160), .A3(new_n1059), .A4(new_n1028), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1056), .A2(new_n1064), .A3(G301), .A4(new_n1057), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1062), .A2(KEYINPUT54), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n959), .A2(G2090), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1971), .B1(new_n967), .B2(new_n969), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(G166), .B2(new_n1034), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1072));
  NAND3_X1  g647(.A1(G303), .A2(G8), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1034), .B1(new_n956), .B2(new_n979), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G305), .A2(G1981), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n574), .A2(new_n1079), .A3(new_n579), .A4(new_n575), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1078), .A2(new_n1080), .A3(new_n1085), .A4(KEYINPUT49), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1077), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n570), .A2(G1976), .A3(new_n571), .A4(new_n572), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n980), .A2(G8), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n996), .A2(G2090), .ZN(new_n1097));
  OAI211_X1 g672(.A(G8), .B(new_n1074), .C1(new_n1097), .C2(new_n1068), .ZN(new_n1098));
  INV_X1    g673(.A(G1976), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1077), .A2(new_n1090), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1076), .A2(new_n1096), .A3(new_n1098), .A4(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT126), .B(KEYINPUT54), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1056), .A2(new_n1057), .A3(new_n1064), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G171), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1056), .A2(G301), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1066), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1024), .A2(new_n1053), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1088), .A2(new_n1099), .A3(new_n760), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1080), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1077), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1098), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1033), .A2(G286), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1102), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1113), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  OAI21_X1  g695(.A(G8), .B1(new_n1097), .B2(new_n1068), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1075), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1119), .A2(new_n1098), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1114), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1109), .A2(KEYINPUT127), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT127), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1105), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1041), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(G168), .A3(new_n1039), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1130), .A2(new_n1046), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT62), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1102), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1048), .A2(new_n1134), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1135));
  AND4_X1   g710(.A1(new_n1127), .A2(new_n1132), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1125), .A2(new_n1126), .A3(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n951), .A2(new_n940), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n586), .B(G1986), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n934), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n955), .B1(new_n1137), .B2(new_n1140), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g716(.A(G319), .ZN(new_n1143));
  OR2_X1    g717(.A1(G229), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g718(.A(new_n1144), .B1(new_n905), .B2(new_n909), .ZN(new_n1145));
  NOR2_X1   g719(.A1(G401), .A2(G227), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n849), .A2(new_n1145), .A3(new_n1146), .ZN(G225));
  INV_X1    g721(.A(G225), .ZN(G308));
endmodule


