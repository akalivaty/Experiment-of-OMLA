//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1235, new_n1236, new_n1237, new_n1238;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT66), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(KEYINPUT66), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n454), .A2(G567), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n478), .B(new_n481), .C1(new_n487), .C2(G124), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n464), .B2(new_n465), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n482), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n492), .B2(new_n494), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT69), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .A3(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(new_n512), .B1(KEYINPUT5), .B2(new_n509), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(G88), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(G50), .A3(G543), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(new_n513), .A2(new_n517), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n529), .A2(G51), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n513), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT74), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(G168));
  NAND2_X1  g117(.A1(new_n510), .A2(new_n512), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(new_n535), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(G64), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n515), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n525), .A2(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n528), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  AOI22_X1  g129(.A1(new_n536), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n515), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n529), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n545), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n570));
  AND2_X1   g145(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n513), .A2(G91), .A3(new_n517), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n573), .A2(new_n576), .ZN(G299));
  XNOR2_X1  g152(.A(G171), .B(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n523), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n516), .B(new_n582), .C1(new_n521), .C2(new_n522), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(G303));
  NAND3_X1  g159(.A1(new_n513), .A2(G87), .A3(new_n517), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(G74), .B1(new_n546), .B2(new_n547), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n587), .B1(new_n589), .B2(G651), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  NAND3_X1  g166(.A1(new_n513), .A2(G86), .A3(new_n517), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n543), .A2(G61), .A3(new_n544), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n598), .A2(new_n599), .A3(G651), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT80), .B1(new_n601), .B2(new_n515), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n594), .A2(new_n595), .A3(new_n600), .A4(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n529), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n515), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(new_n525), .A2(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n545), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n578), .B2(G868), .ZN(G284));
  AOI21_X1  g195(.A(new_n619), .B1(new_n578), .B2(G868), .ZN(G321));
  NOR2_X1   g196(.A1(G299), .A2(G868), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g198(.A(new_n622), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(new_n618), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NOR2_X1   g202(.A1(new_n558), .A2(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n625), .A2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT83), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n631), .B2(G868), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n482), .A2(new_n470), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n487), .A2(G123), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n463), .A2(G111), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(KEYINPUT84), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(KEYINPUT84), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n640), .A2(new_n642), .B1(new_n476), .B2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n637), .A2(G2100), .B1(G2096), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n636), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n645), .B(new_n647), .C1(G2096), .C2(new_n644), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2443), .B(G2446), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT85), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n663), .B(G14), .C1(new_n661), .C2(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n646), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n679), .A2(new_n681), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n684), .A3(new_n682), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n686), .B(new_n689), .C1(new_n684), .C2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT32), .B(G1981), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT90), .B(G16), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n590), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n703), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G24), .B(G290), .S(new_n705), .Z(new_n717));
  INV_X1    g292(.A(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n715), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n487), .A2(G119), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n476), .A2(G131), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n463), .A2(G107), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT88), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n722), .B1(new_n729), .B2(new_n721), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT89), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n730), .B(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n716), .A2(new_n719), .A3(new_n720), .A4(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT92), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n738), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n476), .A2(G139), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n482), .A2(G127), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n463), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n721), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n721), .B2(G33), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n721), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n721), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G2078), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT24), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n721), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G160), .B2(new_n721), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n756), .A2(new_n759), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  NOR2_X1   g345(.A1(G171), .A2(new_n709), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G5), .B2(new_n709), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G4), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n625), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1348), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n772), .A2(new_n770), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n704), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n776), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n784), .A2(new_n721), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n787), .B1(new_n721), .B2(new_n644), .C1(new_n753), .C2(new_n754), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G2078), .B2(new_n758), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n721), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n487), .A2(G128), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n476), .A2(G140), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT94), .ZN(new_n794));
  OR2_X1    g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n791), .B1(new_n798), .B2(new_n721), .ZN(new_n799));
  INV_X1    g374(.A(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n721), .A2(G35), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n721), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT29), .ZN(new_n804));
  INV_X1    g379(.A(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n789), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n704), .A2(G19), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT93), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n559), .B2(new_n704), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1341), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G21), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G168), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1966), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n773), .A2(new_n783), .A3(new_n807), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n721), .A2(G32), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n484), .A2(G129), .A3(new_n486), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n470), .A2(G105), .ZN(new_n822));
  NAND3_X1  g397(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT26), .ZN(new_n824));
  AOI211_X1 g399(.A(new_n822), .B(new_n824), .C1(G141), .C2(new_n476), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n820), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n821), .B1(new_n820), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n817), .B1(new_n828), .B2(new_n721), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT27), .ZN(new_n830));
  INV_X1    g405(.A(G1996), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n816), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n742), .A2(new_n833), .ZN(G311));
  NAND2_X1  g409(.A1(new_n742), .A2(new_n833), .ZN(G150));
  AOI22_X1  g410(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n515), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n525), .A2(G93), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT99), .B(G55), .Z(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n528), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n837), .A2(KEYINPUT100), .A3(new_n840), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT100), .B1(new_n837), .B2(new_n840), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n559), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n559), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT38), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n846), .A2(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n558), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n559), .A2(new_n846), .A3(new_n847), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n618), .A2(new_n626), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n850), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n845), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n861), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n844), .B1(new_n865), .B2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n504), .B(KEYINPUT103), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n826), .B2(new_n827), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n820), .A2(new_n825), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT98), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n820), .A2(new_n821), .A3(new_n825), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n870), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n872), .A2(new_n876), .A3(new_n798), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n798), .B1(new_n872), .B2(new_n876), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n869), .B(new_n751), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n797), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n751), .A2(new_n869), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n750), .A2(KEYINPUT104), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n872), .A2(new_n876), .A3(new_n798), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n487), .A2(G130), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT105), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n476), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n463), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n727), .B(new_n635), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n891), .B(new_n892), .Z(new_n893));
  NAND3_X1  g468(.A1(new_n879), .A2(new_n885), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n879), .B2(new_n885), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n644), .B(G160), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT107), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  INV_X1    g476(.A(new_n899), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n901), .B(new_n902), .C1(new_n895), .C2(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT106), .B(G37), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n897), .B2(new_n899), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n868), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n879), .A2(new_n885), .ZN(new_n910));
  INV_X1    g485(.A(new_n893), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n894), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n901), .B1(new_n913), .B2(new_n902), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n907), .B(new_n868), .C1(new_n909), .C2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n908), .A2(new_n916), .ZN(G395));
  INV_X1    g492(.A(G868), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n842), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G288), .B(G305), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n608), .A2(new_n523), .A3(new_n609), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n523), .B1(new_n608), .B2(new_n609), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n920), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n928), .A2(KEYINPUT109), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n929), .A2(KEYINPUT109), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(KEYINPUT109), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n852), .A2(new_n854), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n630), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n618), .A2(G299), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n618), .A2(G299), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(KEYINPUT41), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n938), .A2(new_n630), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n940), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n943), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n940), .B2(new_n948), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n937), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n934), .B(new_n935), .C1(new_n949), .C2(new_n951), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n936), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n919), .B1(new_n955), .B2(new_n918), .ZN(G295));
  OAI21_X1  g531(.A(new_n919), .B1(new_n955), .B2(new_n918), .ZN(G331));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n578), .A2(G168), .ZN(new_n959));
  OR2_X1    g534(.A1(G168), .A2(G171), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n848), .B2(new_n849), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n852), .A2(new_n854), .A3(new_n959), .A4(new_n960), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n962), .A2(new_n950), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n947), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT112), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT112), .B1(new_n925), .B2(new_n927), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n963), .ZN(new_n970));
  INV_X1    g545(.A(new_n947), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(new_n963), .A3(new_n950), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(KEYINPUT111), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n966), .A2(new_n969), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n964), .A2(new_n965), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n928), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT43), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n964), .A2(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n972), .A2(new_n928), .A3(new_n973), .ZN(new_n980));
  AND4_X1   g555(.A1(KEYINPUT43), .A2(new_n979), .A3(new_n905), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n983), .A2(new_n979), .A3(new_n905), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(new_n977), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(KEYINPUT43), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n986), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g562(.A(KEYINPUT127), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n469), .A2(new_n471), .ZN(new_n989));
  INV_X1    g564(.A(G125), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n474), .B2(new_n475), .ZN(new_n991));
  INV_X1    g566(.A(new_n467), .ZN(new_n992));
  OAI21_X1  g567(.A(G2105), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n993), .A3(G40), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(G160), .A2(KEYINPUT113), .A3(G40), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n504), .B2(G1384), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n797), .B(new_n800), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n828), .B2(new_n831), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n831), .B2(new_n828), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n727), .B(new_n733), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(G290), .B(new_n718), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1001), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  INV_X1    g586(.A(G1971), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n506), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n495), .B2(new_n500), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT45), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(new_n996), .A3(new_n997), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n504), .A2(G1384), .A3(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n495), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1013), .B1(new_n1022), .B2(new_n501), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n996), .A2(new_n997), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n805), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1011), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n581), .A2(G8), .A3(new_n583), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n581), .A2(KEYINPUT55), .A3(G8), .A4(new_n583), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1027), .A2(KEYINPUT115), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT115), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n592), .A2(new_n595), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n602), .A2(new_n600), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G1981), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1981), .B1(new_n529), .B2(G48), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n594), .A2(new_n600), .A3(new_n602), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1040), .A3(KEYINPUT49), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n996), .A2(new_n997), .A3(new_n1015), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT117), .B(KEYINPUT49), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n590), .B2(G1976), .ZN(new_n1052));
  INV_X1    g627(.A(new_n587), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(G1976), .C1(new_n588), .C2(new_n515), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1042), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1050), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G288), .A2(G1976), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1050), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1040), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1035), .A2(new_n1063), .B1(new_n1066), .B2(new_n1043), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  INV_X1    g643(.A(G1966), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT45), .B(new_n1013), .C1(new_n1022), .C2(new_n501), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1025), .A2(new_n1070), .A3(new_n1000), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n998), .A2(G2084), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1069), .A2(new_n1071), .B1(new_n1024), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1011), .B1(new_n1073), .B2(G168), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1069), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1024), .A2(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G286), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1068), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(new_n1076), .A3(G168), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1073), .A2(G168), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT51), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1074), .A2(new_n1068), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1027), .A2(new_n1032), .A3(KEYINPUT115), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G2078), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1025), .A2(new_n1070), .A3(new_n1095), .A4(new_n1000), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1000), .A2(new_n996), .A3(new_n997), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(KEYINPUT123), .A3(new_n1095), .A4(new_n1070), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(KEYINPUT53), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1023), .A2(new_n999), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1016), .A3(new_n1025), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1104), .B2(G2078), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n770), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n578), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n998), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1013), .C1(new_n1022), .C2(new_n501), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1112), .A2(new_n805), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1011), .B1(new_n1018), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1032), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1062), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1094), .A2(new_n1110), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1067), .B1(new_n1089), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G168), .A2(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1073), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1094), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1122), .B(KEYINPUT63), .C1(new_n1032), .C2(new_n1027), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1062), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1123), .A2(new_n1124), .B1(new_n1094), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n573), .B2(new_n576), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT120), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(new_n1129), .C1(new_n573), .C2(new_n576), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1131), .B(new_n1133), .C1(new_n1134), .C2(G299), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1103), .A2(new_n1016), .A3(new_n1025), .A4(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(KEYINPUT118), .B(G1956), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1111), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1025), .A2(new_n1114), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1141), .B2(new_n781), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1135), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n781), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1141), .A2(new_n1139), .A3(new_n781), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT121), .A3(new_n1137), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1135), .B(new_n1137), .C1(new_n1138), .C2(new_n1142), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1042), .A2(G2067), .ZN(new_n1152));
  INV_X1    g727(.A(G1348), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1106), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n618), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1145), .A2(new_n1150), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1135), .B1(new_n1149), .B2(new_n1137), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1151), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n625), .B1(new_n1154), .B2(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1154), .A2(KEYINPUT60), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1154), .A2(KEYINPUT60), .A3(new_n625), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT122), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1042), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1104), .B2(G1996), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1170), .B2(new_n559), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1170), .A2(new_n559), .ZN(new_n1172));
  XNOR2_X1  g747(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1160), .A2(new_n1165), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1151), .A2(KEYINPUT61), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1156), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1101), .A2(G301), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1102), .A2(G2078), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1016), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n994), .B(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1182), .A2(KEYINPUT125), .A3(new_n1184), .A4(new_n1000), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1016), .A2(new_n1000), .A3(new_n1181), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n994), .B(KEYINPUT124), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1190), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1180), .B1(new_n1191), .B2(G171), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1179), .A2(new_n1192), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1193));
  NAND4_X1  g768(.A1(G301), .A2(new_n1190), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1109), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1180), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1050), .B(new_n1061), .C1(new_n1032), .C2(new_n1116), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1193), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1178), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1010), .B1(new_n1128), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1001), .A2(new_n831), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT46), .Z(new_n1203));
  NAND2_X1  g778(.A1(new_n828), .A2(new_n1002), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1203), .B1(new_n1001), .B2(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT47), .Z(new_n1206));
  NAND3_X1  g781(.A1(new_n1004), .A2(new_n729), .A3(new_n733), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(G2067), .B2(new_n797), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1001), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1006), .A2(new_n1001), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n608), .A2(new_n718), .A3(new_n609), .A4(new_n1001), .ZN(new_n1211));
  XOR2_X1   g786(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1212));
  XNOR2_X1  g787(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1206), .A2(new_n1209), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n988), .B1(new_n1201), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1193), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1177), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1218), .A2(new_n1165), .A3(new_n1160), .A4(new_n1174), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1217), .B1(new_n1219), .B2(new_n1156), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1198), .A2(new_n1110), .A3(new_n1083), .A4(new_n1088), .ZN(new_n1221));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n1198), .B2(new_n1122), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1035), .A2(new_n1062), .A3(new_n1125), .ZN(new_n1223));
  OAI211_X1 g798(.A(new_n1221), .B(new_n1067), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1009), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1215), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1225), .A2(KEYINPUT127), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1216), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g803(.A(new_n905), .B1(new_n913), .B2(new_n902), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n1230), .B1(new_n900), .B2(new_n903), .ZN(new_n1231));
  NOR2_X1   g805(.A1(G227), .A2(new_n461), .ZN(new_n1232));
  NAND4_X1  g806(.A1(new_n698), .A2(new_n664), .A3(new_n699), .A4(new_n1232), .ZN(new_n1233));
  NOR3_X1   g807(.A1(new_n986), .A2(new_n1231), .A3(new_n1233), .ZN(G308));
  INV_X1    g808(.A(new_n984), .ZN(new_n1235));
  INV_X1    g809(.A(new_n985), .ZN(new_n1236));
  OAI21_X1  g810(.A(new_n1235), .B1(new_n1236), .B2(new_n983), .ZN(new_n1237));
  NOR2_X1   g811(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1238));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1238), .ZN(G225));
endmodule


