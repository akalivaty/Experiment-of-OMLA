//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n457), .A2(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G101), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G137), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n462), .B(KEYINPUT68), .C1(new_n464), .C2(new_n463), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(G160));
  NOR2_X1   g051(.A1(new_n471), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT70), .Z(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n457), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(G124), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n479), .A2(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n463), .B2(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT71), .A3(new_n489), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n501), .A3(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n495), .A2(new_n497), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT72), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n507), .A2(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n529), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT5), .B(G543), .Z(new_n537));
  NAND2_X1  g112(.A1(new_n512), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G168));
  INV_X1    g118(.A(new_n519), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(G90), .A2(new_n544), .B1(new_n547), .B2(G651), .ZN(new_n548));
  INV_X1    g123(.A(new_n513), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AND2_X1   g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n518), .B2(G56), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n523), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n512), .A2(G43), .A3(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n512), .A2(G81), .A3(new_n518), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(KEYINPUT74), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n554), .C2(new_n523), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n537), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT75), .A3(G651), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n523), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n512), .A2(new_n579), .A3(G53), .A4(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n578), .A2(new_n580), .B1(new_n544), .B2(G91), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G299));
  NAND3_X1  g157(.A1(new_n536), .A2(KEYINPUT76), .A3(new_n541), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n535), .B2(new_n540), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  OAI21_X1  g163(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT77), .Z(new_n590));
  AOI22_X1  g165(.A1(G87), .A2(new_n544), .B1(new_n549), .B2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n516), .B2(new_n517), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n512), .A2(G86), .A3(new_n518), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n544), .A2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n549), .A2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(new_n523), .C2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n537), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(G54), .A2(new_n549), .B1(new_n609), .B2(G651), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n519), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n512), .A2(new_n518), .A3(KEYINPUT10), .A4(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n586), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n586), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n616), .A2(G559), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n625), .A2(KEYINPUT80), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n617), .A2(new_n623), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n562), .A2(new_n626), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n493), .A2(new_n458), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n485), .A2(G123), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G111), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n643), .A2(new_n644), .B1(new_n646), .B2(G2105), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n477), .A2(G135), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n638), .A2(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(G2096), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n639), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT84), .Z(new_n656));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n656), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1341), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1348), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  INV_X1    g254(.A(new_n672), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(new_n691), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n695), .B(new_n697), .C1(new_n687), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT88), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT89), .ZN(new_n702));
  XOR2_X1   g277(.A(G1981), .B(G1986), .Z(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n702), .B(new_n707), .ZN(G229));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT29), .B(G2090), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(G26), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n477), .A2(G140), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G128), .ZN(new_n717));
  OR2_X1    g292(.A1(G104), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G116), .C2(new_n457), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2067), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n713), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT90), .B(G16), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G19), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  INV_X1    g302(.A(new_n725), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n562), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1341), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT23), .Z(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1956), .ZN(new_n734));
  NOR2_X1   g309(.A1(G4), .A2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n616), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1348), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n724), .A2(new_n730), .A3(new_n734), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(G23), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G288), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT33), .B(G1976), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G6), .A2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G305), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT32), .B(G1981), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n743), .ZN(new_n752));
  INV_X1    g327(.A(new_n744), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(new_n748), .B2(new_n749), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n728), .A2(G22), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G166), .B2(new_n728), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1971), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT34), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT34), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n751), .A2(new_n754), .A3(new_n760), .A4(new_n757), .ZN(new_n761));
  MUX2_X1   g336(.A(G24), .B(G290), .S(new_n728), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1986), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n485), .A2(G119), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n457), .A2(G107), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n766));
  INV_X1    g341(.A(G131), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n493), .A2(new_n457), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n764), .B1(new_n765), .B2(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G25), .B(new_n769), .S(G29), .Z(new_n770));
  XOR2_X1   g345(.A(KEYINPUT35), .B(G1991), .Z(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n770), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n763), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n759), .A2(new_n761), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n775), .A2(KEYINPUT91), .A3(KEYINPUT36), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n759), .A2(new_n777), .A3(new_n761), .A4(new_n774), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n740), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT102), .ZN(new_n780));
  OR2_X1    g355(.A1(G29), .A2(G33), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n457), .A2(G103), .A3(G2104), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n768), .ZN(new_n786));
  NAND2_X1  g361(.A1(G115), .A2(G2104), .ZN(new_n787));
  INV_X1    g362(.A(G127), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n471), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n786), .B1(G2105), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT95), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n790), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n781), .B1(new_n797), .B2(new_n709), .ZN(new_n798));
  INV_X1    g373(.A(G2072), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n737), .A2(G21), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n542), .B2(G16), .ZN(new_n801));
  INV_X1    g376(.A(G1966), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n798), .A2(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n709), .A2(G32), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n458), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n485), .A2(G129), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT26), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n807), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT27), .B(G1996), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n801), .A2(new_n802), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n737), .A2(G5), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G301), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(G1961), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n709), .A2(G27), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G164), .B2(new_n709), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G2078), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(G2078), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n823), .A2(new_n824), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n825), .A2(new_n828), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n816), .A2(new_n818), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT30), .B(G28), .ZN(new_n833));
  OR2_X1    g408(.A1(KEYINPUT31), .A2(G11), .ZN(new_n834));
  NAND2_X1  g409(.A1(KEYINPUT31), .A2(G11), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n833), .A2(new_n709), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n649), .B2(new_n709), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR4_X1   g414(.A1(new_n821), .A2(new_n831), .A3(new_n832), .A4(new_n839), .ZN(new_n840));
  OAI211_X1 g415(.A(G2072), .B(new_n781), .C1(new_n797), .C2(new_n709), .ZN(new_n841));
  OR2_X1    g416(.A1(KEYINPUT24), .A2(G34), .ZN(new_n842));
  NAND2_X1  g417(.A1(KEYINPUT24), .A2(G34), .ZN(new_n843));
  AOI21_X1  g418(.A(G29), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G160), .B2(G29), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(G2084), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n806), .A2(new_n840), .A3(new_n841), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(G2084), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n780), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n806), .A2(new_n841), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(KEYINPUT97), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n840), .A2(new_n848), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(KEYINPUT102), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n779), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(G311));
  XNOR2_X1  g434(.A(new_n858), .B(KEYINPUT103), .ZN(G150));
  XNOR2_X1  g435(.A(KEYINPUT105), .B(G55), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n549), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G67), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n516), .B2(new_n517), .ZN(new_n864));
  AND2_X1   g439(.A1(G80), .A2(G543), .ZN(new_n865));
  OAI21_X1  g440(.A(G651), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n512), .A2(G93), .A3(new_n518), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n558), .A2(new_n561), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n862), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n559), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n617), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g453(.A(G860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n870), .A2(G860), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT37), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(G145));
  XNOR2_X1  g458(.A(G160), .B(new_n649), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(G162), .Z(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n813), .A2(new_n814), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(new_n720), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n815), .A2(new_n721), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n505), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n888), .A2(new_n505), .A3(new_n889), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n792), .B(new_n796), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n769), .B(new_n636), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n485), .A2(G130), .ZN(new_n895));
  OR2_X1    g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(G2104), .C1(G118), .C2(new_n457), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G142), .B2(new_n477), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n894), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n892), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n794), .A3(new_n890), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n893), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n893), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n886), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n891), .A2(new_n791), .A3(new_n892), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n797), .B1(new_n902), .B2(new_n890), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n900), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n904), .A3(new_n885), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(G303), .A2(G305), .ZN(new_n915));
  NAND2_X1  g490(.A1(G166), .A2(new_n747), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(KEYINPUT110), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(KEYINPUT110), .A3(new_n916), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G288), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n918), .B(new_n919), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n924), .A2(new_n923), .A3(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n576), .A2(new_n581), .A3(new_n610), .A4(new_n615), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n576), .A2(new_n581), .B1(new_n610), .B2(new_n615), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT41), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g508(.A1(G299), .A2(new_n616), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n929), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n562), .A2(new_n870), .ZN(new_n938));
  INV_X1    g513(.A(new_n871), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n629), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n625), .B1(new_n869), .B2(new_n871), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n930), .A2(new_n931), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(KEYINPUT107), .A3(new_n935), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n937), .A2(new_n942), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n937), .A2(new_n942), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n928), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n947), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT42), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n927), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n928), .A3(new_n950), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT42), .B1(new_n952), .B2(new_n953), .ZN(new_n957));
  INV_X1    g532(.A(new_n927), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n626), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n870), .A2(new_n626), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n960), .A2(KEYINPUT111), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n958), .B1(new_n956), .B2(new_n957), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n961), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(G295));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n961), .ZN(G331));
  AOI21_X1  g545(.A(G301), .B1(new_n583), .B2(new_n585), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n541), .A2(new_n536), .B1(new_n548), .B2(new_n550), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n938), .A2(new_n939), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n872), .B1(new_n971), .B2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n943), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n937), .A2(new_n944), .A3(new_n975), .A4(new_n976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT112), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n975), .A2(new_n976), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n944), .A4(new_n937), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n958), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n977), .B1(new_n936), .B2(new_n932), .ZN(new_n987));
  INV_X1    g562(.A(new_n978), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n927), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n985), .A2(new_n986), .A3(new_n908), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT113), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n984), .B2(new_n958), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n986), .A4(new_n989), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n980), .A2(new_n927), .A3(new_n983), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n985), .A2(new_n908), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n992), .A2(KEYINPUT43), .A3(new_n989), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT43), .B1(new_n992), .B2(new_n995), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(G397));
  AOI21_X1  g579(.A(KEYINPUT71), .B1(new_n493), .B2(new_n489), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n503), .B1(new_n496), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1006), .B2(new_n495), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT45), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n468), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT68), .B1(new_n493), .B2(new_n462), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n459), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n470), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n493), .B2(G125), .ZN(new_n1014));
  OAI21_X1  g589(.A(G40), .B1(new_n1014), .B2(new_n457), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G40), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n473), .B2(G2105), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n469), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1009), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1996), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n887), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2067), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n720), .B(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n815), .A2(G1996), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n769), .A2(new_n772), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n769), .A2(new_n772), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G290), .B(G1986), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1022), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n598), .A2(new_n1036), .A3(new_n599), .A4(new_n600), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT116), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1035), .A2(new_n1041), .A3(KEYINPUT49), .A4(new_n1037), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1007), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(G8), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G288), .A2(G1976), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1046), .A2(new_n1047), .B1(new_n1036), .B2(new_n747), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n922), .A2(G1976), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(new_n1052), .A3(G8), .A4(new_n1044), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(new_n1051), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1046), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G1384), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n505), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(new_n1021), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1018), .A2(new_n469), .A3(new_n1019), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1019), .B1(new_n1018), .B2(new_n469), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1384), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n497), .A2(new_n502), .A3(new_n498), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT50), .ZN(new_n1073));
  NOR2_X1   g648(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1065), .A2(G1971), .B1(new_n1076), .B2(G2090), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1060), .A2(new_n1077), .A3(G8), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1048), .A2(new_n1049), .B1(new_n1056), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(KEYINPUT63), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1046), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(G8), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1059), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1084), .A3(new_n1078), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1072), .A2(new_n1061), .B1(new_n505), .B2(new_n1062), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1966), .B1(new_n1086), .B2(new_n1068), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1075), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n505), .B2(new_n1069), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1088), .A2(G2084), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G286), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1081), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1056), .B1(new_n1083), .B2(new_n1059), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1081), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(new_n1078), .A3(new_n1097), .A4(new_n1093), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1079), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n802), .B1(new_n1064), .B2(new_n1021), .ZN(new_n1101));
  INV_X1    g676(.A(G2084), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1068), .A2(new_n1102), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n542), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1101), .A2(new_n1104), .A3(new_n1103), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1104), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1113));
  OAI21_X1  g688(.A(G168), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1109), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1092), .B(new_n1107), .C1(new_n1108), .C2(G168), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G168), .A2(new_n1108), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1100), .A2(new_n1119), .A3(new_n1105), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G2078), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT53), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1012), .A2(new_n1015), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1009), .A2(KEYINPUT125), .A3(new_n1063), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1063), .A2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1008), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1086), .A2(new_n1068), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(G2078), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n824), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n1134), .B2(KEYINPUT126), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(KEYINPUT126), .B2(new_n1134), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1132), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1133), .B1(new_n1131), .B2(new_n1123), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1133), .B(new_n1141), .C1(new_n1131), .C2(new_n1123), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1137), .B1(new_n1143), .B2(G301), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1136), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1129), .A2(new_n1132), .A3(G301), .A4(new_n1133), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1143), .B2(G301), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1085), .B1(new_n1147), .B2(new_n1137), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1121), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n576), .B2(new_n581), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1086), .A2(new_n1068), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G1956), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1348), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1068), .A2(new_n1025), .A3(new_n1007), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n616), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1153), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT118), .B(G1996), .Z(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1086), .A2(new_n1068), .A3(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1044), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n563), .A3(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(KEYINPUT120), .B(new_n562), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1173), .A2(new_n563), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(KEYINPUT120), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT121), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1158), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1153), .B1(new_n1157), .B2(new_n1155), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1166), .A2(new_n1158), .A3(KEYINPUT61), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1160), .A2(new_n616), .A3(new_n1161), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT60), .B1(new_n1188), .B2(new_n1162), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1160), .A2(new_n1161), .A3(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1182), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1178), .A2(KEYINPUT121), .A3(new_n1181), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1167), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1099), .B1(new_n1149), .B2(new_n1195), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1085), .A2(G301), .A3(new_n1143), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1121), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1118), .A2(KEYINPUT62), .A3(new_n1120), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1034), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(G290), .A2(G1986), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1022), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT48), .Z(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n1032), .B2(new_n1022), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT46), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1026), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1022), .B1(new_n815), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT47), .Z(new_n1212));
  OAI22_X1  g787(.A1(new_n1028), .A2(new_n1031), .B1(G2067), .B2(new_n720), .ZN(new_n1213));
  AOI211_X1 g788(.A(new_n1206), .B(new_n1212), .C1(new_n1022), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1202), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g790(.A1(new_n684), .A2(G319), .ZN(new_n1217));
  XOR2_X1   g791(.A(new_n1217), .B(KEYINPUT127), .Z(new_n1218));
  NOR3_X1   g792(.A1(G229), .A2(G401), .A3(new_n1218), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n998), .A2(new_n1219), .A3(new_n913), .ZN(G308));
  NAND3_X1  g794(.A1(new_n998), .A2(new_n1219), .A3(new_n913), .ZN(G225));
endmodule


