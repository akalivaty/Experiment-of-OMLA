

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748;

  XNOR2_X1 U370 ( .A(n373), .B(n372), .ZN(n408) );
  OR2_X1 U371 ( .A1(n544), .A2(n682), .ZN(n529) );
  AND2_X1 U372 ( .A1(n418), .A2(n527), .ZN(n349) );
  XNOR2_X1 U373 ( .A(n737), .B(n432), .ZN(n503) );
  XNOR2_X1 U374 ( .A(n402), .B(G119), .ZN(n497) );
  XNOR2_X1 U375 ( .A(n442), .B(n428), .ZN(n514) );
  INV_X2 U376 ( .A(G953), .ZN(n739) );
  XNOR2_X2 U377 ( .A(n576), .B(KEYINPUT66), .ZN(n577) );
  NAND2_X2 U378 ( .A1(n378), .A2(n377), .ZN(n658) );
  NAND2_X1 U379 ( .A1(n349), .A2(n590), .ZN(n544) );
  NAND2_X1 U380 ( .A1(n583), .A2(n581), .ZN(n582) );
  XNOR2_X2 U381 ( .A(n578), .B(n577), .ZN(n583) );
  XOR2_X1 U382 ( .A(n555), .B(KEYINPUT43), .Z(n350) );
  AND2_X2 U383 ( .A1(n393), .A2(n395), .ZN(n392) );
  XNOR2_X2 U384 ( .A(n505), .B(n427), .ZN(n722) );
  XNOR2_X2 U385 ( .A(n497), .B(n496), .ZN(n505) );
  NOR2_X1 U386 ( .A1(n560), .A2(n666), .ZN(n587) );
  AND2_X1 U387 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U388 ( .A1(n379), .A2(KEYINPUT85), .ZN(n377) );
  AND2_X1 U389 ( .A1(n624), .A2(n638), .ZN(n585) );
  OR2_X1 U390 ( .A1(n380), .A2(n534), .ZN(n382) );
  NOR2_X1 U391 ( .A1(n547), .A2(n540), .ZN(n639) );
  NAND2_X1 U392 ( .A1(n547), .A2(n540), .ZN(n647) );
  AND2_X1 U393 ( .A1(n595), .A2(n403), .ZN(n531) );
  XNOR2_X1 U394 ( .A(n457), .B(n456), .ZN(n547) );
  XNOR2_X1 U395 ( .A(n405), .B(n491), .ZN(n595) );
  XOR2_X1 U396 ( .A(n703), .B(KEYINPUT59), .Z(n704) );
  XNOR2_X1 U397 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  INV_X1 U398 ( .A(KEYINPUT89), .ZN(n495) );
  XNOR2_X1 U399 ( .A(n582), .B(KEYINPUT32), .ZN(n351) );
  NAND2_X1 U400 ( .A1(n705), .A2(n704), .ZN(n354) );
  NAND2_X1 U401 ( .A1(n352), .A2(n353), .ZN(n355) );
  NAND2_X1 U402 ( .A1(n354), .A2(n355), .ZN(n706) );
  INV_X1 U403 ( .A(n705), .ZN(n352) );
  INV_X1 U404 ( .A(n704), .ZN(n353) );
  BUF_X1 U405 ( .A(n714), .Z(n356) );
  XNOR2_X1 U406 ( .A(n582), .B(KEYINPUT32), .ZN(n624) );
  NOR2_X1 U407 ( .A1(n706), .A2(n720), .ZN(n709) );
  NAND2_X1 U408 ( .A1(n383), .A2(n360), .ZN(n578) );
  NAND2_X1 U409 ( .A1(n386), .A2(n384), .ZN(n426) );
  NAND2_X1 U410 ( .A1(n387), .A2(n645), .ZN(n386) );
  XNOR2_X1 U411 ( .A(n538), .B(n362), .ZN(n422) );
  XNOR2_X1 U412 ( .A(n514), .B(n431), .ZN(n737) );
  XNOR2_X1 U413 ( .A(n430), .B(n429), .ZN(n431) );
  INV_X1 U414 ( .A(G137), .ZN(n429) );
  XNOR2_X1 U415 ( .A(G131), .B(G134), .ZN(n430) );
  XNOR2_X1 U416 ( .A(n409), .B(n441), .ZN(n534) );
  XNOR2_X1 U417 ( .A(n421), .B(n420), .ZN(n379) );
  NOR2_X1 U418 ( .A1(n426), .A2(n424), .ZN(n423) );
  OR2_X1 U419 ( .A1(n746), .A2(KEYINPUT85), .ZN(n375) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n498) );
  XOR2_X1 U421 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n446) );
  XNOR2_X1 U422 ( .A(KEYINPUT105), .B(KEYINPUT7), .ZN(n445) );
  XOR2_X1 U423 ( .A(KEYINPUT103), .B(G122), .Z(n444) );
  NAND2_X1 U424 ( .A1(n532), .A2(n525), .ZN(n419) );
  XNOR2_X1 U425 ( .A(n433), .B(n411), .ZN(n721) );
  XNOR2_X1 U426 ( .A(G104), .B(G107), .ZN(n433) );
  XNOR2_X1 U427 ( .A(n412), .B(G110), .ZN(n411) );
  INV_X1 U428 ( .A(KEYINPUT77), .ZN(n412) );
  XNOR2_X1 U429 ( .A(KEYINPUT79), .B(KEYINPUT88), .ZN(n509) );
  XNOR2_X1 U430 ( .A(n721), .B(n410), .ZN(n437) );
  INV_X1 U431 ( .A(KEYINPUT73), .ZN(n410) );
  XNOR2_X1 U432 ( .A(n374), .B(n363), .ZN(n696) );
  AND2_X1 U433 ( .A1(n389), .A2(n596), .ZN(n553) );
  NOR2_X1 U434 ( .A1(n647), .A2(n390), .ZN(n389) );
  INV_X1 U435 ( .A(n531), .ZN(n390) );
  XNOR2_X1 U436 ( .A(n534), .B(KEYINPUT1), .ZN(n560) );
  INV_X1 U437 ( .A(KEYINPUT28), .ZN(n381) );
  INV_X1 U438 ( .A(n592), .ZN(n672) );
  NAND2_X2 U439 ( .A1(n392), .A2(n391), .ZN(n383) );
  NAND2_X1 U440 ( .A1(n370), .A2(n357), .ZN(n391) );
  XNOR2_X1 U441 ( .A(n592), .B(KEYINPUT6), .ZN(n596) );
  NOR2_X1 U442 ( .A1(n551), .A2(KEYINPUT47), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n550), .B(n425), .ZN(n424) );
  INV_X1 U444 ( .A(KEYINPUT81), .ZN(n425) );
  INV_X1 U445 ( .A(G237), .ZN(n515) );
  AND2_X1 U446 ( .A1(n376), .A2(n361), .ZN(n378) );
  XOR2_X1 U447 ( .A(KEYINPUT12), .B(G122), .Z(n459) );
  XNOR2_X1 U448 ( .A(G113), .B(G131), .ZN(n458) );
  XOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n462) );
  XNOR2_X1 U450 ( .A(G143), .B(G104), .ZN(n464) );
  XNOR2_X1 U451 ( .A(n506), .B(n406), .ZN(n485) );
  XNOR2_X1 U452 ( .A(G140), .B(KEYINPUT10), .ZN(n406) );
  XOR2_X1 U453 ( .A(KEYINPUT70), .B(G101), .Z(n507) );
  XNOR2_X1 U454 ( .A(n407), .B(G125), .ZN(n506) );
  INV_X1 U455 ( .A(G146), .ZN(n407) );
  NAND2_X1 U456 ( .A1(G234), .A2(G237), .ZN(n470) );
  INV_X1 U457 ( .A(n668), .ZN(n404) );
  INV_X1 U458 ( .A(n570), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n503), .B(n502), .ZN(n610) );
  XNOR2_X1 U460 ( .A(n500), .B(n499), .ZN(n501) );
  BUF_X1 U461 ( .A(n658), .Z(n738) );
  XNOR2_X1 U462 ( .A(G116), .B(G107), .ZN(n443) );
  INV_X1 U463 ( .A(n560), .ZN(n579) );
  XNOR2_X1 U464 ( .A(n419), .B(n364), .ZN(n418) );
  INV_X1 U465 ( .A(n595), .ZN(n669) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n626) );
  XNOR2_X1 U467 ( .A(n437), .B(n512), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n722), .B(n400), .ZN(n399) );
  INV_X1 U469 ( .A(n382), .ZN(n539) );
  NOR2_X1 U470 ( .A1(n385), .A2(n560), .ZN(n652) );
  XNOR2_X1 U471 ( .A(n524), .B(KEYINPUT36), .ZN(n385) );
  INV_X1 U472 ( .A(KEYINPUT35), .ZN(n372) );
  INV_X1 U473 ( .A(n676), .ZN(n416) );
  AND2_X1 U474 ( .A1(n394), .A2(n572), .ZN(n357) );
  NOR2_X1 U475 ( .A1(n547), .A2(n546), .ZN(n358) );
  AND2_X1 U476 ( .A1(n746), .A2(KEYINPUT85), .ZN(n359) );
  AND2_X1 U477 ( .A1(n683), .A2(n668), .ZN(n360) );
  AND2_X1 U478 ( .A1(n375), .A2(n655), .ZN(n361) );
  XNOR2_X1 U479 ( .A(KEYINPUT64), .B(n537), .ZN(n362) );
  XOR2_X1 U480 ( .A(n564), .B(n563), .Z(n363) );
  XNOR2_X1 U481 ( .A(KEYINPUT30), .B(KEYINPUT113), .ZN(n364) );
  XNOR2_X1 U482 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n365) );
  NOR2_X1 U483 ( .A1(n739), .A2(G952), .ZN(n720) );
  XNOR2_X1 U484 ( .A(n413), .B(n365), .ZN(n366) );
  XNOR2_X1 U485 ( .A(n413), .B(n365), .ZN(n396) );
  NAND2_X1 U486 ( .A1(n367), .A2(n608), .ZN(n609) );
  NAND2_X1 U487 ( .A1(n368), .A2(n605), .ZN(n367) );
  NAND2_X1 U488 ( .A1(n396), .A2(n369), .ZN(n368) );
  NOR2_X1 U489 ( .A1(n658), .A2(n602), .ZN(n369) );
  NAND2_X1 U490 ( .A1(n371), .A2(n417), .ZN(n393) );
  INV_X1 U491 ( .A(n371), .ZN(n370) );
  NOR2_X1 U492 ( .A1(n371), .A2(n382), .ZN(n645) );
  XNOR2_X2 U493 ( .A(n397), .B(KEYINPUT19), .ZN(n371) );
  NAND2_X1 U494 ( .A1(n626), .A2(n602), .ZN(n520) );
  NAND2_X1 U495 ( .A1(n575), .A2(n358), .ZN(n373) );
  NAND2_X1 U496 ( .A1(n562), .A2(n596), .ZN(n374) );
  NOR2_X1 U497 ( .A1(n616), .A2(G902), .ZN(n409) );
  NAND2_X1 U498 ( .A1(n379), .A2(n359), .ZN(n376) );
  XNOR2_X1 U499 ( .A(n533), .B(n381), .ZN(n380) );
  XNOR2_X2 U500 ( .A(n523), .B(KEYINPUT87), .ZN(n397) );
  NAND2_X1 U501 ( .A1(n383), .A2(n590), .ZN(n591) );
  NAND2_X1 U502 ( .A1(n383), .A2(n416), .ZN(n589) );
  NAND2_X1 U503 ( .A1(n696), .A2(n383), .ZN(n574) );
  INV_X1 U504 ( .A(n652), .ZN(n384) );
  XNOR2_X1 U505 ( .A(n388), .B(KEYINPUT76), .ZN(n387) );
  NAND2_X1 U506 ( .A1(n570), .A2(n417), .ZN(n395) );
  INV_X1 U507 ( .A(n366), .ZN(n726) );
  NAND2_X1 U508 ( .A1(n607), .A2(n366), .ZN(n608) );
  NAND2_X1 U509 ( .A1(n553), .A2(n397), .ZN(n524) );
  XNOR2_X1 U510 ( .A(n401), .B(n513), .ZN(n400) );
  INV_X1 U511 ( .A(n514), .ZN(n401) );
  XNOR2_X2 U512 ( .A(G116), .B(KEYINPUT3), .ZN(n402) );
  NOR2_X1 U513 ( .A1(n526), .A2(n404), .ZN(n403) );
  NOR2_X1 U514 ( .A1(n716), .A2(G902), .ZN(n405) );
  NAND2_X1 U515 ( .A1(n585), .A2(n408), .ZN(n415) );
  XNOR2_X1 U516 ( .A(n408), .B(G122), .ZN(G24) );
  NAND2_X2 U517 ( .A1(n414), .A2(n601), .ZN(n413) );
  XNOR2_X2 U518 ( .A(n415), .B(n586), .ZN(n414) );
  INV_X1 U519 ( .A(n572), .ZN(n417) );
  XNOR2_X2 U520 ( .A(n504), .B(G472), .ZN(n532) );
  INV_X1 U521 ( .A(KEYINPUT48), .ZN(n420) );
  NAND2_X1 U522 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U523 ( .A(n620), .B(n619), .ZN(n622) );
  XNOR2_X1 U524 ( .A(n503), .B(n438), .ZN(n616) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(G122), .Z(n427) );
  INV_X1 U526 ( .A(KEYINPUT5), .ZN(n499) );
  INV_X1 U527 ( .A(KEYINPUT109), .ZN(n561) );
  XNOR2_X1 U528 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U529 ( .A(G469), .ZN(n439) );
  XNOR2_X1 U530 ( .A(n480), .B(n481), .ZN(n484) );
  XNOR2_X1 U531 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U532 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U533 ( .A(G146), .B(n507), .ZN(n432) );
  XOR2_X2 U534 ( .A(G143), .B(G128), .Z(n442) );
  INV_X1 U535 ( .A(KEYINPUT4), .ZN(n428) );
  XOR2_X1 U536 ( .A(G140), .B(KEYINPUT78), .Z(n435) );
  NAND2_X1 U537 ( .A1(G227), .A2(n739), .ZN(n434) );
  XNOR2_X1 U538 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U540 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n440) );
  XNOR2_X1 U541 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n455) );
  XNOR2_X1 U542 ( .A(n442), .B(G134), .ZN(n453) );
  XNOR2_X1 U543 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U544 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U545 ( .A(n448), .B(n447), .Z(n451) );
  NAND2_X1 U546 ( .A1(G234), .A2(n739), .ZN(n449) );
  XOR2_X1 U547 ( .A(KEYINPUT8), .B(n449), .Z(n482) );
  NAND2_X1 U548 ( .A1(G217), .A2(n482), .ZN(n450) );
  XNOR2_X1 U549 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U550 ( .A(n453), .B(n452), .ZN(n710) );
  NOR2_X1 U551 ( .A1(G902), .A2(n710), .ZN(n454) );
  XNOR2_X1 U552 ( .A(n455), .B(n454), .ZN(n457) );
  INV_X1 U553 ( .A(G478), .ZN(n456) );
  XNOR2_X1 U554 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U555 ( .A(n485), .B(n460), .ZN(n467) );
  NAND2_X1 U556 ( .A1(G214), .A2(n498), .ZN(n461) );
  XNOR2_X1 U557 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U558 ( .A(n463), .B(KEYINPUT101), .Z(n465) );
  XNOR2_X1 U559 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U560 ( .A(n467), .B(n466), .ZN(n703) );
  NOR2_X1 U561 ( .A1(G902), .A2(n703), .ZN(n469) );
  XOR2_X1 U562 ( .A(KEYINPUT13), .B(G475), .Z(n468) );
  XNOR2_X1 U563 ( .A(n469), .B(n468), .ZN(n546) );
  INV_X1 U564 ( .A(n546), .ZN(n540) );
  XNOR2_X1 U565 ( .A(n470), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U566 ( .A1(G952), .A2(n473), .ZN(n694) );
  NOR2_X1 U567 ( .A1(G953), .A2(n694), .ZN(n472) );
  INV_X1 U568 ( .A(KEYINPUT92), .ZN(n471) );
  XNOR2_X1 U569 ( .A(n472), .B(n471), .ZN(n569) );
  INV_X1 U570 ( .A(n569), .ZN(n477) );
  NAND2_X1 U571 ( .A1(n473), .A2(G902), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n474), .B(KEYINPUT95), .ZN(n566) );
  NAND2_X1 U573 ( .A1(n566), .A2(G953), .ZN(n475) );
  NOR2_X1 U574 ( .A1(G900), .A2(n475), .ZN(n476) );
  NOR2_X1 U575 ( .A1(n477), .A2(n476), .ZN(n526) );
  XOR2_X1 U576 ( .A(G110), .B(G128), .Z(n481) );
  XOR2_X1 U577 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n479) );
  XNOR2_X1 U578 ( .A(G119), .B(G137), .ZN(n478) );
  NAND2_X1 U579 ( .A1(G221), .A2(n482), .ZN(n483) );
  XNOR2_X1 U580 ( .A(n484), .B(n483), .ZN(n486) );
  INV_X1 U581 ( .A(n485), .ZN(n736) );
  XNOR2_X1 U582 ( .A(n486), .B(n736), .ZN(n716) );
  NAND2_X1 U583 ( .A1(n602), .A2(G234), .ZN(n488) );
  XNOR2_X1 U584 ( .A(KEYINPUT20), .B(KEYINPUT98), .ZN(n487) );
  XNOR2_X1 U585 ( .A(n488), .B(n487), .ZN(n492) );
  NAND2_X1 U586 ( .A1(G217), .A2(n492), .ZN(n490) );
  XNOR2_X1 U587 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n489) );
  XNOR2_X1 U588 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U589 ( .A1(n492), .A2(G221), .ZN(n494) );
  INV_X1 U590 ( .A(KEYINPUT21), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n494), .B(n493), .ZN(n668) );
  XNOR2_X1 U592 ( .A(n495), .B(G113), .ZN(n496) );
  NAND2_X1 U593 ( .A1(n498), .A2(G210), .ZN(n500) );
  XNOR2_X1 U594 ( .A(n505), .B(n501), .ZN(n502) );
  INV_X1 U595 ( .A(G902), .ZN(n516) );
  NAND2_X1 U596 ( .A1(n610), .A2(n516), .ZN(n504) );
  INV_X1 U597 ( .A(n532), .ZN(n592) );
  XNOR2_X1 U598 ( .A(n507), .B(n506), .ZN(n513) );
  NAND2_X1 U599 ( .A1(n739), .A2(G224), .ZN(n508) );
  XNOR2_X1 U600 ( .A(n509), .B(n508), .ZN(n511) );
  XNOR2_X1 U601 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n510) );
  XNOR2_X1 U602 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U603 ( .A1(n516), .A2(n515), .ZN(n521) );
  NAND2_X1 U604 ( .A1(n521), .A2(G210), .ZN(n518) );
  INV_X1 U605 ( .A(KEYINPUT90), .ZN(n517) );
  XNOR2_X1 U606 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X2 U607 ( .A(n520), .B(n519), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n521), .A2(G214), .ZN(n522) );
  XNOR2_X1 U609 ( .A(n522), .B(KEYINPUT91), .ZN(n681) );
  INV_X1 U610 ( .A(n681), .ZN(n525) );
  NAND2_X1 U611 ( .A1(n543), .A2(n525), .ZN(n523) );
  NAND2_X1 U612 ( .A1(n669), .A2(n668), .ZN(n666) );
  NOR2_X1 U613 ( .A1(n534), .A2(n666), .ZN(n590) );
  INV_X1 U614 ( .A(n526), .ZN(n527) );
  XNOR2_X1 U615 ( .A(n543), .B(KEYINPUT38), .ZN(n682) );
  XNOR2_X2 U616 ( .A(n529), .B(KEYINPUT39), .ZN(n559) );
  INV_X1 U617 ( .A(n647), .ZN(n644) );
  NAND2_X1 U618 ( .A1(n559), .A2(n644), .ZN(n530) );
  XNOR2_X1 U619 ( .A(n530), .B(KEYINPUT40), .ZN(n747) );
  AND2_X1 U620 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U621 ( .A1(n547), .A2(n546), .ZN(n683) );
  NOR2_X1 U622 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U623 ( .A1(n683), .A2(n686), .ZN(n535) );
  XNOR2_X1 U624 ( .A(n535), .B(KEYINPUT41), .ZN(n695) );
  NAND2_X1 U625 ( .A1(n539), .A2(n695), .ZN(n536) );
  XNOR2_X1 U626 ( .A(n536), .B(KEYINPUT42), .ZN(n748) );
  NAND2_X1 U627 ( .A1(n747), .A2(n748), .ZN(n538) );
  XOR2_X1 U628 ( .A(KEYINPUT46), .B(KEYINPUT86), .Z(n537) );
  XNOR2_X1 U629 ( .A(KEYINPUT108), .B(n639), .ZN(n558) );
  INV_X1 U630 ( .A(n558), .ZN(n541) );
  NAND2_X1 U631 ( .A1(n541), .A2(n647), .ZN(n685) );
  NAND2_X1 U632 ( .A1(n645), .A2(n685), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n542), .A2(KEYINPUT47), .ZN(n549) );
  INV_X1 U634 ( .A(n543), .ZN(n556) );
  NOR2_X1 U635 ( .A1(n544), .A2(n556), .ZN(n545) );
  XNOR2_X1 U636 ( .A(n545), .B(KEYINPUT114), .ZN(n548) );
  NAND2_X1 U637 ( .A1(n548), .A2(n358), .ZN(n642) );
  NAND2_X1 U638 ( .A1(n549), .A2(n642), .ZN(n550) );
  INV_X1 U639 ( .A(n685), .ZN(n551) );
  NOR2_X1 U640 ( .A1(n681), .A2(n579), .ZN(n552) );
  NAND2_X1 U641 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U642 ( .A(KEYINPUT111), .B(n554), .ZN(n555) );
  NAND2_X1 U643 ( .A1(n350), .A2(n556), .ZN(n557) );
  XNOR2_X1 U644 ( .A(n557), .B(KEYINPUT112), .ZN(n746) );
  NAND2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n655) );
  XNOR2_X1 U646 ( .A(n587), .B(n561), .ZN(n562) );
  XNOR2_X1 U647 ( .A(KEYINPUT110), .B(KEYINPUT33), .ZN(n564) );
  INV_X1 U648 ( .A(KEYINPUT74), .ZN(n563) );
  XNOR2_X1 U649 ( .A(G898), .B(KEYINPUT93), .ZN(n729) );
  NAND2_X1 U650 ( .A1(n729), .A2(G953), .ZN(n565) );
  XOR2_X1 U651 ( .A(KEYINPUT94), .B(n565), .Z(n724) );
  NAND2_X1 U652 ( .A1(n566), .A2(n724), .ZN(n567) );
  XNOR2_X1 U653 ( .A(n567), .B(KEYINPUT96), .ZN(n568) );
  AND2_X1 U654 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U655 ( .A(KEYINPUT69), .ZN(n571) );
  XNOR2_X1 U656 ( .A(n571), .B(KEYINPUT0), .ZN(n572) );
  INV_X1 U657 ( .A(KEYINPUT34), .ZN(n573) );
  XNOR2_X1 U658 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n576) );
  NAND2_X1 U660 ( .A1(n579), .A2(n595), .ZN(n580) );
  NOR2_X1 U661 ( .A1(n580), .A2(n596), .ZN(n581) );
  AND2_X1 U662 ( .A1(n583), .A2(n560), .ZN(n598) );
  NOR2_X1 U663 ( .A1(n672), .A2(n669), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n598), .A2(n584), .ZN(n638) );
  INV_X1 U665 ( .A(KEYINPUT44), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n672), .ZN(n676) );
  XOR2_X1 U667 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n588) );
  XNOR2_X1 U668 ( .A(n589), .B(n588), .ZN(n650) );
  XNOR2_X1 U669 ( .A(n591), .B(KEYINPUT99), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n634) );
  NAND2_X1 U671 ( .A1(n650), .A2(n634), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n594), .A2(n685), .ZN(n600) );
  NOR2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  AND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n631) );
  INV_X1 U675 ( .A(n631), .ZN(n599) );
  AND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT83), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  XOR2_X1 U679 ( .A(KEYINPUT67), .B(n604), .Z(n605) );
  INV_X1 U680 ( .A(KEYINPUT2), .ZN(n606) );
  NOR2_X1 U681 ( .A1(n658), .A2(n606), .ZN(n607) );
  XNOR2_X2 U682 ( .A(n609), .B(KEYINPUT65), .ZN(n714) );
  NAND2_X1 U683 ( .A1(n714), .A2(G472), .ZN(n612) );
  XOR2_X1 U684 ( .A(KEYINPUT62), .B(n610), .Z(n611) );
  XNOR2_X1 U685 ( .A(n612), .B(n611), .ZN(n613) );
  INV_X1 U686 ( .A(n613), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(n621), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U689 ( .A1(n714), .A2(G469), .ZN(n620) );
  XOR2_X1 U690 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n618) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT121), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n619) );
  INV_X1 U693 ( .A(n720), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT122), .ZN(G54) );
  XNOR2_X1 U695 ( .A(n351), .B(G119), .ZN(G21) );
  NAND2_X1 U696 ( .A1(n714), .A2(G210), .ZN(n628) );
  XNOR2_X1 U697 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X2 U700 ( .A1(n629), .A2(n720), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U702 ( .A(G101), .B(n631), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT115), .ZN(G3) );
  NOR2_X1 U704 ( .A1(n647), .A2(n634), .ZN(n633) );
  XOR2_X1 U705 ( .A(G104), .B(n633), .Z(G6) );
  INV_X1 U706 ( .A(n639), .ZN(n649) );
  NOR2_X1 U707 ( .A1(n649), .A2(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U710 ( .A(G107), .B(n637), .ZN(G9) );
  XNOR2_X1 U711 ( .A(n638), .B(G110), .ZN(G12) );
  XOR2_X1 U712 ( .A(G128), .B(KEYINPUT29), .Z(n641) );
  NAND2_X1 U713 ( .A1(n645), .A2(n639), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G30) );
  XNOR2_X1 U715 ( .A(G143), .B(KEYINPUT116), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(G45) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(G146), .B(n646), .ZN(G48) );
  NOR2_X1 U719 ( .A1(n650), .A2(n647), .ZN(n648) );
  XOR2_X1 U720 ( .A(G113), .B(n648), .Z(G15) );
  NOR2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(G116), .B(n651), .Z(G18) );
  XOR2_X1 U723 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n654) );
  XNOR2_X1 U724 ( .A(G125), .B(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(G27) );
  XNOR2_X1 U726 ( .A(G134), .B(n655), .ZN(G36) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n656) );
  NAND2_X1 U728 ( .A1(n726), .A2(n656), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT82), .ZN(n664) );
  NAND2_X1 U730 ( .A1(KEYINPUT80), .A2(n738), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT2), .ZN(n662) );
  INV_X1 U732 ( .A(n738), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n660), .A2(n726), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n665), .A2(n739), .ZN(n701) );
  NAND2_X1 U737 ( .A1(n666), .A2(n560), .ZN(n667) );
  XNOR2_X1 U738 ( .A(KEYINPUT50), .B(n667), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(n670), .Z(n671) );
  NOR2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n675), .B(KEYINPUT118), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U745 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n695), .A2(n680), .ZN(n691) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n696), .A2(n689), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U754 ( .A(KEYINPUT52), .B(n692), .Z(n693) );
  NOR2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n698) );
  AND2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U758 ( .A(KEYINPUT120), .B(n699), .Z(n700) );
  NOR2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U760 ( .A(KEYINPUT53), .B(n702), .ZN(G75) );
  NAND2_X1 U761 ( .A1(n714), .A2(G475), .ZN(n705) );
  XOR2_X1 U762 ( .A(KEYINPUT60), .B(KEYINPUT68), .Z(n707) );
  XNOR2_X1 U763 ( .A(KEYINPUT123), .B(n707), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(G60) );
  NAND2_X1 U765 ( .A1(n356), .A2(G478), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n710), .B(KEYINPUT124), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n720), .A2(n713), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n356), .A2(G217), .ZN(n718) );
  INV_X1 U770 ( .A(KEYINPUT125), .ZN(n715) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n720), .A2(n719), .ZN(G66) );
  XOR2_X1 U773 ( .A(n721), .B(G101), .Z(n723) );
  XNOR2_X1 U774 ( .A(n722), .B(n723), .ZN(n725) );
  NOR2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n734) );
  NOR2_X1 U776 ( .A1(n726), .A2(G953), .ZN(n732) );
  XOR2_X1 U777 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n728) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n730) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U781 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U782 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U783 ( .A(KEYINPUT127), .B(n735), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n741), .B(n738), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n745) );
  XNOR2_X1 U787 ( .A(G227), .B(n741), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(G953), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n745), .A2(n744), .ZN(G72) );
  XNOR2_X1 U791 ( .A(G140), .B(n746), .ZN(G42) );
  XNOR2_X1 U792 ( .A(n747), .B(G131), .ZN(G33) );
  XNOR2_X1 U793 ( .A(G137), .B(n748), .ZN(G39) );
endmodule

