//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AND2_X1   g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G97), .A2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n202), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n211), .B(new_n214), .C1(G87), .C2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G50), .A2(G226), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n225), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n226), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n248), .A2(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n226), .B1(new_n201), .B2(new_n203), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n247), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n226), .A2(G1), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n247), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n255), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G222), .B2(G1698), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G77), .B2(new_n274), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G226), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n276), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G200), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT10), .B1(new_n268), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n265), .A2(new_n289), .A3(new_n266), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT10), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n284), .B(new_n292), .C1(new_n285), .C2(new_n283), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT68), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n296), .B(new_n293), .C1(new_n288), .C2(new_n290), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n287), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G97), .ZN(new_n299));
  INV_X1    g0099(.A(G226), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G232), .B2(new_n301), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n299), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n270), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n278), .A2(G238), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n282), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G200), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n317), .B(KEYINPUT69), .Z(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n313), .A2(new_n319), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G190), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n249), .A2(new_n202), .B1(new_n226), .B2(G68), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT71), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n259), .B2(new_n252), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n247), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n326), .B2(new_n247), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n330), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(KEYINPUT11), .A3(new_n328), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT66), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n261), .A2(new_n334), .A3(G13), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n337), .A2(new_n261), .A3(new_n247), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT12), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(KEYINPUT12), .A3(new_n220), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n257), .A2(new_n339), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AND4_X1   g0143(.A1(new_n322), .A2(new_n331), .A3(new_n333), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n331), .A2(new_n333), .A3(new_n343), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n315), .A2(G169), .A3(new_n316), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT14), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n320), .A2(G179), .A3(new_n321), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n315), .A2(new_n349), .A3(G169), .A4(new_n316), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n318), .A2(new_n344), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n283), .A2(G179), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n283), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n263), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G20), .A2(G77), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT15), .B(G87), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n357), .B1(new_n252), .B2(new_n248), .C1(new_n359), .C2(new_n249), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n247), .B1(new_n338), .B2(G77), .ZN(new_n361));
  INV_X1    g0161(.A(new_n337), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(G77), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n221), .A2(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G232), .B2(G1698), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n270), .B1(new_n365), .B2(new_n274), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G107), .B2(new_n274), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n278), .A2(G244), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n282), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n354), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n363), .B(new_n370), .C1(G179), .C2(new_n369), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n298), .A2(new_n352), .A3(new_n356), .A4(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT7), .B1(new_n274), .B2(G20), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n308), .A2(new_n374), .A3(new_n226), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n375), .A3(G68), .ZN(new_n376));
  XNOR2_X1  g0176(.A(G58), .B(G68), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n304), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n307), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT75), .B1(new_n304), .B2(KEYINPUT3), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT7), .B(new_n226), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n374), .B1(new_n274), .B2(G20), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n220), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n378), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n376), .A2(KEYINPUT74), .A3(KEYINPUT16), .A4(new_n378), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n381), .A2(new_n390), .A3(new_n247), .A4(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n248), .A2(new_n247), .A3(new_n261), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n258), .B2(new_n248), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n271), .A2(new_n301), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n300), .A2(G1698), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n305), .A2(new_n396), .A3(new_n307), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n310), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT76), .ZN(new_n402));
  INV_X1    g0202(.A(G179), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n281), .B1(new_n278), .B2(G232), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n405), .A3(new_n310), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n354), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n395), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n395), .A2(new_n411), .A3(KEYINPUT18), .ZN(new_n415));
  INV_X1    g0215(.A(G200), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(G190), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n392), .A2(new_n419), .A3(new_n394), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n392), .A2(new_n419), .A3(new_n394), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT77), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n414), .A2(new_n415), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n369), .A2(G200), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n369), .A2(new_n285), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n363), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n372), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G97), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G107), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(KEYINPUT6), .B1(new_n435), .B2(G107), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT6), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT78), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n435), .A2(G107), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n439), .A2(KEYINPUT6), .ZN(new_n445));
  AND4_X1   g0245(.A1(new_n438), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n437), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n445), .ZN(new_n448));
  INV_X1    g0248(.A(new_n442), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT79), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n440), .A2(new_n438), .A3(new_n442), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(new_n436), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n447), .A2(G20), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n251), .A2(G77), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n386), .A2(new_n387), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G107), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n247), .ZN(new_n458));
  INV_X1    g0258(.A(new_n247), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n256), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n257), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n462), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G97), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n258), .A2(new_n435), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n458), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(new_n301), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n310), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  INV_X1    g0277(.A(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(G274), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n225), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n477), .A2(new_n479), .B1(new_n481), .B2(new_n269), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G257), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n484), .A2(G179), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n354), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n468), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n457), .A2(new_n247), .B1(G97), .B2(new_n465), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(G200), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n476), .A2(G190), .A3(new_n480), .A4(new_n483), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n467), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n274), .A2(new_n226), .A3(G68), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT19), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n249), .B2(new_n435), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n226), .B1(new_n299), .B2(new_n493), .ZN(new_n497));
  INV_X1    g0297(.A(G87), .ZN(new_n498));
  INV_X1    g0298(.A(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n435), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n497), .A2(KEYINPUT82), .A3(new_n500), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n495), .A2(new_n496), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n503), .A2(new_n492), .A3(new_n494), .A4(new_n504), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n507), .A3(new_n247), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n465), .A2(new_n358), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n337), .A2(new_n359), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n221), .A2(new_n301), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n213), .A2(G1698), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n274), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n270), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n479), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n280), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(G250), .A3(new_n270), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n403), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n354), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n511), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR4_X1   g0325(.A1(new_n516), .A2(new_n520), .A3(new_n285), .A4(new_n518), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(G200), .B2(new_n521), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n465), .A2(G87), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n510), .A3(new_n508), .A4(new_n528), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n487), .A2(new_n491), .A3(new_n525), .A4(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n531), .A2(new_n226), .A3(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT23), .B1(new_n499), .B2(G20), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n305), .A2(new_n307), .A3(new_n226), .A4(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n274), .A2(new_n537), .A3(new_n226), .A4(G87), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(KEYINPUT24), .A3(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n247), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n499), .B1(new_n463), .B2(new_n464), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n258), .B(new_n499), .C1(new_n548), .C2(KEYINPUT88), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(KEYINPUT88), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n305), .A2(new_n307), .A3(G250), .A4(new_n301), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n305), .A2(new_n307), .A3(G257), .A4(G1698), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n554), .C1(new_n304), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n310), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT89), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n482), .B2(G264), .ZN(new_n559));
  INV_X1    g0359(.A(G41), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT5), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT5), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G41), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n479), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G264), .A3(new_n270), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(KEYINPUT89), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n557), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT90), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n557), .B(KEYINPUT90), .C1(new_n559), .C2(new_n566), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n480), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n416), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n557), .B(new_n480), .C1(new_n559), .C2(new_n566), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n552), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n536), .A2(new_n538), .ZN(new_n577));
  INV_X1    g0377(.A(new_n534), .ZN(new_n578));
  AND4_X1   g0378(.A1(KEYINPUT24), .A2(new_n577), .A3(new_n540), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT24), .B1(new_n539), .B2(new_n540), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n546), .B1(new_n581), .B2(new_n247), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n569), .A2(G179), .A3(new_n480), .A4(new_n570), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n573), .A2(G169), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(new_n551), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT91), .B1(new_n576), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n552), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT91), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n574), .B1(new_n571), .B2(new_n416), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n589), .C1(new_n552), .C2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n305), .A2(new_n307), .A3(G264), .A4(G1698), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT84), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n274), .A2(new_n594), .A3(G264), .A4(G1698), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n274), .A2(G257), .A3(new_n301), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n308), .A2(G303), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n310), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n482), .A2(G270), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n480), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n362), .A2(G116), .A3(new_n459), .A4(new_n460), .ZN(new_n602));
  INV_X1    g0402(.A(G116), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n246), .A2(new_n225), .B1(G20), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n473), .B(new_n226), .C1(G33), .C2(new_n435), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n606), .A2(KEYINPUT20), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(KEYINPUT20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n604), .A2(new_n606), .A3(new_n605), .A4(KEYINPUT20), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT85), .B1(new_n337), .B2(new_n603), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n337), .A2(KEYINPUT85), .A3(new_n603), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n602), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n601), .A2(new_n615), .A3(G169), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n601), .A2(new_n403), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n615), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n601), .A2(new_n615), .A3(KEYINPUT21), .A4(G169), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n615), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n601), .A2(new_n285), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(G200), .B2(new_n601), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n530), .A2(new_n586), .A3(new_n591), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n434), .A2(new_n627), .ZN(G372));
  NAND2_X1  g0428(.A1(new_n414), .A2(new_n415), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n351), .A2(new_n345), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n371), .B1(new_n422), .B2(new_n427), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n318), .A2(new_n344), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n298), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n356), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n622), .A2(KEYINPUT92), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n618), .A2(new_n620), .A3(new_n639), .A4(new_n621), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n588), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n576), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n641), .A2(new_n530), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n525), .A2(new_n529), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n468), .A2(new_n485), .A3(new_n486), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT26), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n525), .A2(new_n529), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n647), .A2(new_n487), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n525), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n637), .B1(new_n434), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT93), .ZN(G369));
  INV_X1    g0453(.A(G13), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n256), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n626), .B1(new_n623), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n638), .A2(new_n640), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n623), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT94), .B(G330), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n552), .A2(new_n661), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n586), .A2(new_n591), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n585), .A2(new_n661), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT95), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT95), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n670), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n588), .A2(new_n661), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n622), .A2(KEYINPUT96), .A3(new_n662), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT96), .B1(new_n622), .B2(new_n662), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n674), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n208), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G1), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n500), .A2(G116), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n228), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n695), .B(new_n662), .C1(new_n643), .C2(new_n650), .ZN(new_n696));
  INV_X1    g0496(.A(new_n525), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT26), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n648), .B1(new_n647), .B2(new_n487), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n585), .A2(new_n622), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n530), .A2(new_n701), .A3(new_n642), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n661), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n696), .B1(new_n695), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n484), .A2(new_n403), .A3(new_n601), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n569), .A2(new_n570), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n522), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n522), .A4(new_n706), .ZN(new_n710));
  INV_X1    g0510(.A(new_n571), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n484), .A2(new_n403), .A3(new_n601), .A4(new_n521), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n661), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT31), .B(new_n714), .C1(new_n627), .C2(new_n661), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n716), .A3(new_n661), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n704), .B1(new_n668), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n694), .B1(new_n719), .B2(G1), .ZN(G364));
  OR2_X1    g0520(.A1(new_n667), .A2(new_n668), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n691), .B1(G45), .B2(new_n655), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n669), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT97), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n229), .A2(new_n478), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n688), .A2(new_n274), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(new_n244), .C2(new_n478), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n274), .A2(G355), .A3(new_n208), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(G116), .C2(new_n208), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n225), .B1(G20), .B2(new_n354), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT98), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n226), .A2(new_n285), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n403), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n226), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G322), .A2(new_n741), .B1(new_n745), .B2(G329), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n226), .B1(new_n743), .B2(G190), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n746), .B(new_n308), .C1(new_n555), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n403), .A2(new_n416), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n742), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n739), .A2(new_n742), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(new_n752), .B1(new_n754), .B2(G311), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n416), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n742), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n738), .A2(new_n749), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n755), .B1(new_n756), .B2(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n738), .A2(new_n757), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n748), .B(new_n761), .C1(G303), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n745), .A2(G159), .ZN(new_n765));
  INV_X1    g0565(.A(new_n760), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n765), .A2(KEYINPUT32), .B1(G50), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n762), .A2(new_n498), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n754), .A2(G77), .ZN(new_n770));
  INV_X1    g0570(.A(new_n747), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G97), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n767), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G58), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n740), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n765), .A2(KEYINPUT32), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n274), .B1(new_n758), .B2(new_n499), .C1(new_n220), .C2(new_n750), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n773), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n732), .B1(new_n764), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n735), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n737), .B(new_n779), .C1(new_n667), .C2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n725), .B1(new_n723), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT99), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n718), .A2(new_n668), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n641), .A2(new_n530), .A3(new_n642), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n661), .B1(new_n785), .B2(new_n700), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n371), .A2(new_n661), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n363), .A2(new_n661), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n431), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n789), .B2(new_n371), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n786), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n723), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT102), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n784), .A2(new_n792), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(KEYINPUT102), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n791), .A2(new_n734), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n756), .A2(new_n750), .B1(new_n740), .B2(new_n555), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n772), .A2(new_n308), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G303), .C2(new_n766), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n763), .A2(G107), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n758), .A2(new_n498), .B1(new_n744), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT100), .Z(new_n805));
  NAND2_X1  g0605(.A1(new_n754), .A2(G116), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n801), .A2(new_n802), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G143), .A2(new_n741), .B1(new_n754), .B2(G159), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n809), .B2(new_n760), .C1(new_n250), .C2(new_n750), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G58), .B2(new_n771), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n758), .A2(new_n220), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n745), .A2(G132), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n763), .A2(G50), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n807), .B1(new_n817), .B2(new_n308), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n732), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n732), .A2(new_n733), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n202), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n798), .A2(new_n722), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n797), .A2(new_n822), .ZN(G384));
  INV_X1    g0623(.A(new_n659), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n395), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n428), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n412), .A2(new_n825), .A3(new_n423), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n412), .A2(new_n825), .A3(new_n829), .A4(new_n423), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT38), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n376), .A2(new_n378), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n382), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n381), .A2(new_n834), .A3(new_n247), .A4(new_n391), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n394), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n428), .A2(new_n659), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n392), .A2(new_n419), .A3(new_n394), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n835), .A2(new_n394), .B1(new_n410), .B2(new_n659), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT104), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT104), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(KEYINPUT37), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(new_n830), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT105), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT105), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n842), .A2(new_n847), .A3(new_n830), .A4(new_n844), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n838), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n832), .B1(new_n849), .B2(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n345), .A2(new_n661), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n352), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n351), .A2(new_n345), .A3(new_n661), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n715), .A2(new_n717), .A3(new_n854), .A4(new_n791), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT40), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND4_X1   g0657(.A1(new_n715), .A2(new_n717), .A3(new_n791), .A4(new_n854), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n859), .B(new_n838), .C1(new_n846), .C2(new_n848), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n846), .A2(new_n848), .ZN(new_n861));
  INV_X1    g0661(.A(new_n838), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n858), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n857), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n718), .A2(new_n433), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n668), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n631), .A2(new_n661), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT39), .B1(new_n860), .B2(new_n863), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n850), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n860), .A2(new_n863), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n787), .B1(new_n786), .B2(new_n791), .ZN(new_n878));
  INV_X1    g0678(.A(new_n854), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n877), .A2(new_n880), .B1(new_n630), .B2(new_n659), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n636), .B1(new_n704), .B2(new_n433), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n882), .B(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(KEYINPUT106), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(KEYINPUT106), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n887), .B1(new_n256), .B2(new_n655), .C1(new_n886), .C2(new_n868), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n447), .A2(new_n452), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT35), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n226), .B(new_n225), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(G116), .C1(new_n890), .C2(new_n889), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT36), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n202), .B(new_n228), .C1(G58), .C2(G68), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n201), .A2(G68), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n654), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n893), .B1(new_n256), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n888), .A2(new_n898), .ZN(G367));
  NAND2_X1  g0699(.A1(new_n468), .A2(new_n661), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n487), .A2(new_n491), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT108), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT108), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n487), .A2(new_n900), .A3(new_n903), .A4(new_n491), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n645), .A2(new_n661), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n676), .B2(new_n678), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n674), .A2(new_n685), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n588), .B1(new_n902), .B2(new_n904), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n662), .B1(new_n912), .B2(new_n645), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n508), .A2(new_n510), .A3(new_n528), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n661), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n644), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n525), .B2(new_n915), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n697), .A2(KEYINPUT107), .A3(new_n914), .A4(new_n661), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n911), .A2(new_n913), .B1(KEYINPUT43), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n920), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT43), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n911), .A2(new_n923), .A3(new_n922), .A4(new_n913), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n907), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT110), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n907), .A3(new_n926), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT109), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n689), .B(KEYINPUT41), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n686), .A2(new_n908), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT112), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT112), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n686), .A2(new_n936), .A3(new_n908), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n933), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n686), .B2(new_n908), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n684), .B1(new_n672), .B2(new_n673), .ZN(new_n940));
  NOR4_X1   g0740(.A1(new_n940), .A2(new_n906), .A3(KEYINPUT112), .A4(new_n681), .ZN(new_n941));
  INV_X1    g0741(.A(new_n933), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n906), .B1(new_n940), .B2(new_n681), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(KEYINPUT44), .B(new_n906), .C1(new_n940), .C2(new_n681), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(KEYINPUT113), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT113), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n950), .A3(new_n946), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n679), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n952), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n935), .A2(new_n937), .A3(new_n933), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n942), .B1(new_n939), .B2(new_n941), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n957), .A3(new_n680), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n675), .A2(new_n959), .A3(new_n684), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n684), .B1(new_n675), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n719), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n953), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n932), .B1(new_n965), .B2(new_n719), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n256), .B1(new_n655), .B2(G45), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n928), .B(new_n930), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n723), .B1(new_n922), .B2(new_n735), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n762), .A2(new_n603), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT46), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n274), .B(new_n972), .C1(G283), .C2(new_n754), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n758), .A2(new_n435), .B1(new_n744), .B2(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n760), .A2(new_n803), .B1(new_n750), .B2(new_n555), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(G303), .C2(new_n741), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n973), .B(new_n977), .C1(new_n499), .C2(new_n747), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n274), .B1(new_n744), .B2(new_n809), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n774), .A2(new_n762), .B1(new_n740), .B2(new_n250), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(G68), .C2(new_n771), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n766), .A2(G143), .ZN(new_n982));
  INV_X1    g0782(.A(G159), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n750), .A2(new_n983), .B1(new_n753), .B2(new_n201), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT114), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n758), .A2(new_n202), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(new_n985), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n981), .A2(new_n982), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n978), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n732), .ZN(new_n992));
  INV_X1    g0792(.A(new_n727), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n736), .B1(new_n208), .B2(new_n359), .C1(new_n237), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n970), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n969), .A2(new_n995), .ZN(G387));
  OAI21_X1  g0796(.A(new_n274), .B1(new_n753), .B2(new_n220), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n771), .A2(new_n358), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n259), .B2(new_n740), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n762), .A2(new_n202), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n750), .A2(new_n248), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n758), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n997), .B(new_n1002), .C1(G97), .C2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n250), .B2(new_n744), .C1(new_n983), .C2(new_n760), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G322), .A2(new_n766), .B1(new_n751), .B2(G311), .ZN(new_n1006));
  INV_X1    g0806(.A(G303), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n753), .C1(new_n974), .C2(new_n740), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT48), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n756), .B2(new_n747), .C1(new_n555), .C2(new_n762), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT49), .Z(new_n1011));
  OAI221_X1 g0811(.A(new_n308), .B1(new_n744), .B2(new_n759), .C1(new_n603), .C2(new_n758), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1005), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n732), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n672), .A2(new_n673), .A3(new_n735), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n727), .B1(new_n234), .B2(new_n478), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n692), .A2(new_n208), .A3(new_n274), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n692), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n248), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n208), .A2(G107), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n736), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1014), .A2(new_n1015), .A3(new_n722), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n962), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n689), .B1(new_n1025), .B2(new_n719), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1024), .B1(new_n967), .B2(new_n962), .C1(new_n1026), .C2(new_n964), .ZN(G393));
  NAND3_X1  g0827(.A1(new_n953), .A2(new_n968), .A3(new_n958), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n750), .A2(new_n201), .B1(new_n753), .B2(new_n248), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G77), .B2(new_n771), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT115), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n760), .A2(new_n250), .B1(new_n740), .B2(new_n983), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT51), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n762), .A2(new_n220), .B1(new_n758), .B2(new_n498), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n308), .B(new_n1034), .C1(G143), .C2(new_n745), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n750), .A2(new_n1007), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n760), .A2(new_n974), .B1(new_n740), .B2(new_n803), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n274), .B1(new_n1003), .B2(G107), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n754), .A2(G294), .ZN(new_n1041));
  INV_X1    g0841(.A(G322), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n762), .A2(new_n756), .B1(new_n744), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G116), .B2(new_n771), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1036), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n732), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n736), .B1(new_n435), .B2(new_n208), .C1(new_n241), .C2(new_n993), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n722), .A3(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT116), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n780), .B2(new_n908), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1028), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT117), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1028), .A2(KEYINPUT117), .A3(new_n1051), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n964), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n944), .A2(new_n679), .A3(new_n952), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n680), .B1(new_n954), .B2(new_n957), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT118), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1057), .B(KEYINPUT118), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1062), .A2(new_n689), .A3(new_n965), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1056), .A2(new_n1064), .ZN(G390));
  OAI21_X1  g0865(.A(new_n870), .B1(new_n878), .B2(new_n879), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n871), .A2(new_n873), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n849), .A2(KEYINPUT38), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n832), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n787), .B1(new_n703), .B2(new_n791), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n870), .C1(new_n879), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n715), .A2(new_n668), .A3(new_n717), .A4(new_n791), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n879), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n858), .A2(G330), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n715), .A2(G330), .A3(new_n717), .A4(new_n791), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(new_n879), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(new_n1075), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1074), .A2(new_n879), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n878), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1071), .A2(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(KEYINPUT29), .B(new_n661), .C1(new_n785), .C2(new_n700), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n700), .A2(new_n702), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n695), .B1(new_n1087), .B2(new_n662), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n433), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n433), .A2(G330), .A3(new_n715), .A4(new_n717), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n637), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT119), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n883), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1076), .A2(new_n1078), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1077), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1073), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1093), .B1(new_n883), .B2(new_n1090), .ZN(new_n1099));
  AND4_X1   g0899(.A1(new_n1093), .A2(new_n1089), .A3(new_n1090), .A4(new_n637), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1067), .B(new_n1072), .C1(new_n879), .C2(new_n1074), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1079), .A2(new_n879), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n1071), .C1(new_n879), .C2(new_n1074), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n858), .A2(G330), .B1(new_n1074), .B2(new_n879), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n878), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1096), .A2(new_n689), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1098), .A2(new_n968), .A3(new_n1102), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n871), .A2(new_n733), .A3(new_n873), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n762), .A2(new_n250), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n274), .C1(new_n809), .C2(new_n750), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI22_X1  g0914(.A1(G132), .A2(new_n741), .B1(new_n754), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n983), .B2(new_n747), .C1(new_n201), .C2(new_n758), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n760), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n744), .A2(new_n1119), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1113), .A2(new_n1116), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n766), .A2(G283), .B1(new_n771), .B2(G77), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n435), .B2(new_n753), .C1(new_n603), .C2(new_n740), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n308), .B1(new_n744), .B2(new_n555), .C1(new_n499), .C2(new_n750), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1123), .A2(new_n768), .A3(new_n813), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n732), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n820), .A2(new_n248), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1110), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1108), .B(new_n1109), .C1(new_n723), .C2(new_n1128), .ZN(G378));
  INV_X1    g0929(.A(new_n880), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1130), .A2(new_n876), .B1(new_n629), .B2(new_n824), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n865), .B(G330), .C1(new_n874), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n356), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n635), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n263), .A2(new_n824), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1070), .A2(KEYINPUT40), .A3(new_n858), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n863), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n855), .B1(new_n1140), .B2(new_n1068), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(G330), .C1(new_n1141), .C2(KEYINPUT40), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n875), .A3(new_n881), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1132), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1138), .B1(new_n1132), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n968), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n723), .B1(new_n1138), .B2(new_n733), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n760), .A2(new_n1119), .B1(new_n747), .B2(new_n250), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G132), .A2(new_n751), .B1(new_n754), .B2(G137), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1117), .B2(new_n740), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(new_n763), .C2(new_n1114), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(G41), .B1(new_n745), .B2(G124), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G33), .B1(new_n1003), .B2(G159), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(G50), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n751), .A2(G97), .B1(new_n754), .B2(new_n358), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1003), .A2(G58), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1159), .A2(new_n560), .A3(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n760), .A2(new_n603), .B1(new_n744), .B2(new_n756), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n308), .B1(new_n747), .B2(new_n220), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1162), .A2(new_n1000), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1161), .B(new_n1164), .C1(new_n499), .C2(new_n740), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT58), .Z(new_n1166));
  OAI21_X1  g0966(.A(new_n732), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n820), .A2(new_n201), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1147), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1146), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1138), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1142), .A2(new_n875), .A3(new_n881), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1142), .B1(new_n875), .B2(new_n881), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1132), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1175), .A2(new_n1176), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n689), .B1(new_n1177), .B2(KEYINPUT57), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1107), .A2(new_n1101), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(KEYINPUT57), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1171), .B1(new_n1178), .B2(new_n1181), .ZN(G375));
  NAND2_X1  g0982(.A1(new_n820), .A2(new_n220), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n854), .B2(new_n734), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n998), .B1(new_n435), .B2(new_n762), .C1(new_n1007), .C2(new_n744), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n987), .B(new_n1185), .C1(G283), .C2(new_n741), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n766), .A2(G294), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n754), .A2(G107), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n274), .B1(new_n751), .B2(G116), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n274), .B1(new_n747), .B2(new_n259), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1160), .B1(new_n1117), .B2(new_n744), .C1(new_n983), .C2(new_n762), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G150), .C2(new_n754), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT121), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n766), .A2(G132), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n751), .A2(new_n1114), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n740), .A2(new_n809), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1190), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n723), .B(new_n1184), .C1(new_n732), .C2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1106), .B2(new_n968), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1085), .A2(new_n1095), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n931), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1085), .A2(new_n1095), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(G381));
  OAI21_X1  g1005(.A(new_n1179), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n690), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1170), .B1(new_n1208), .B2(new_n1180), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1109), .B1(new_n723), .B2(new_n1128), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1107), .A2(new_n689), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1096), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1213), .A2(G396), .A3(G393), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n969), .A2(new_n1056), .A3(new_n1064), .A4(new_n995), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(G384), .A3(G381), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n660), .A2(G213), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT122), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(new_n1213), .C2(new_n1219), .ZN(G409));
  NAND2_X1  g1020(.A1(G387), .A2(G390), .ZN(new_n1221));
  XOR2_X1   g1021(.A(G393), .B(G396), .Z(new_n1222));
  AND3_X1   g1022(.A1(new_n1221), .A2(new_n1215), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1221), .B2(new_n1215), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1179), .B(new_n931), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n1212), .A2(new_n1146), .A3(new_n1169), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G375), .B2(G378), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT124), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1202), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n690), .B1(new_n1232), .B2(KEYINPUT60), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1201), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(G384), .A3(new_n1201), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(KEYINPUT125), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1238), .A2(G384), .A3(new_n1201), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1238), .B2(new_n1201), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1228), .A2(new_n1218), .A3(new_n1243), .A4(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT62), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1171), .A2(new_n1212), .A3(new_n1226), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1219), .C1(new_n1209), .C2(new_n1212), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1247), .A2(new_n1243), .A3(KEYINPUT62), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1248), .A2(new_n1249), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n660), .A2(G213), .A3(G2897), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1247), .A2(new_n1243), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1219), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(G2897), .A3(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1225), .B1(new_n1254), .B2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1250), .B(new_n1218), .C1(new_n1209), .C2(new_n1212), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT63), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1248), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1247), .A2(new_n1243), .A3(KEYINPUT63), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1261), .B1(new_n1251), .B2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n1225), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(G405));
  AOI211_X1 g1072(.A(G378), .B(new_n1170), .C1(new_n1208), .C2(new_n1180), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n689), .A3(new_n1180), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1212), .B1(new_n1275), .B2(new_n1171), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1257), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1276), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1280), .A2(new_n1213), .A3(new_n1243), .A4(new_n1247), .ZN(new_n1281));
  OAI211_X1 g1081(.A(KEYINPUT126), .B(new_n1257), .C1(new_n1273), .C2(new_n1276), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1223), .A2(new_n1224), .A3(KEYINPUT127), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1222), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1215), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n995), .A2(new_n969), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1221), .A2(new_n1215), .A3(new_n1222), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1285), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1284), .A2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1283), .B(new_n1292), .ZN(G402));
endmodule


