//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n209), .C1(new_n202), .C2(KEYINPUT1), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT68), .B1(KEYINPUT67), .B2(KEYINPUT28), .ZN(new_n217));
  OR2_X1    g016(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n218));
  AND4_X1   g017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT26), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n220), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n217), .B1(new_n216), .B2(new_n215), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n219), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G183gat), .B(G190gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n230), .B(new_n232), .C1(new_n233), .C2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n222), .B1(new_n220), .B2(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n237), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n215), .A2(G183gat), .ZN(new_n241));
  INV_X1    g040(.A(G183gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G190gat), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT24), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n230), .B1(new_n244), .B2(new_n232), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n229), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n237), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n222), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n231), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n242), .A2(G190gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n215), .A2(G183gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n256), .B2(KEYINPUT24), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n252), .B1(new_n229), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n246), .A2(new_n247), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n247), .B1(new_n246), .B2(new_n258), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n214), .B(new_n228), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n257), .A2(new_n230), .B1(new_n235), .B2(new_n250), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n233), .A2(new_n231), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT64), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT25), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n258), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT66), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n246), .A2(new_n247), .A3(new_n258), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n214), .A4(new_n228), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n228), .B1(new_n259), .B2(new_n260), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n213), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n263), .A2(new_n272), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT32), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n272), .A3(new_n274), .ZN(new_n280));
  INV_X1    g079(.A(new_n275), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT33), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n278), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT33), .B1(new_n280), .B2(new_n281), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n290), .A2(new_n282), .A3(new_n285), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n280), .A2(new_n281), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n286), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n278), .B1(new_n297), .B2(new_n288), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT36), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT2), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n302));
  XNOR2_X1  g101(.A(G155gat), .B(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n301), .ZN(new_n304));
  XNOR2_X1  g103(.A(G141gat), .B(G148gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G141gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G148gat), .ZN(new_n308));
  INV_X1    g107(.A(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n301), .B(new_n311), .C1(new_n314), .C2(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n213), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT5), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n315), .A3(KEYINPUT3), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n322), .A2(new_n213), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n324), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  AOI211_X1 g125(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n306), .C2(new_n315), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n316), .A2(new_n211), .A3(new_n212), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n214), .A2(KEYINPUT4), .A3(new_n316), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n328), .A2(new_n318), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n213), .A2(new_n315), .A3(new_n306), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n329), .ZN(new_n335));
  INV_X1    g134(.A(new_n318), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n328), .A2(new_n341), .A3(new_n318), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n316), .A2(new_n211), .A3(new_n212), .A4(new_n330), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n214), .B2(new_n316), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n340), .B1(new_n342), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n328), .A2(new_n341), .A3(new_n318), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n214), .A2(KEYINPUT81), .A3(new_n316), .A4(new_n330), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n346), .B2(new_n349), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT82), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n339), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G1gat), .B(G29gat), .Z(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT82), .B1(new_n353), .B2(new_n355), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n351), .A3(new_n340), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT79), .B1(new_n337), .B2(KEYINPUT5), .ZN(new_n368));
  AOI211_X1 g167(.A(new_n320), .B(new_n341), .C1(new_n335), .C2(new_n336), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n366), .A2(new_n367), .B1(new_n370), .B2(new_n333), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n365), .B1(new_n371), .B2(new_n362), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n364), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(G211gat), .A2(G218gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G197gat), .B(G204gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT71), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT71), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n377), .C1(new_n380), .C2(new_n381), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT73), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT74), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n227), .B1(new_n269), .B2(new_n270), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n227), .B1(new_n246), .B2(new_n258), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n392), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n273), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n390), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n394), .B1(new_n398), .B2(KEYINPUT29), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n401), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n409), .B(KEYINPUT75), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n392), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n402), .B1(new_n273), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n416), .B2(new_n399), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT30), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n418), .A3(new_n409), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n374), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT31), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G50gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G228gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n325), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n434));
  INV_X1    g233(.A(new_n316), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n326), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n316), .A2(new_n324), .A3(new_n325), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(new_n392), .ZN(new_n440));
  INV_X1    g239(.A(new_n382), .ZN(new_n441));
  INV_X1    g240(.A(new_n386), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n415), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n316), .B1(new_n443), .B2(new_n325), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n415), .B1(new_n326), .B2(new_n327), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n390), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n446), .B2(new_n432), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(G22gat), .ZN(new_n448));
  INV_X1    g247(.A(G22gat), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n440), .B(new_n449), .C1(new_n432), .C2(new_n446), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n425), .B(new_n429), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n450), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n428), .B1(new_n452), .B2(KEYINPUT83), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n425), .A3(new_n450), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n424), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n278), .ZN(new_n458));
  INV_X1    g257(.A(new_n288), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n291), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n297), .A2(new_n278), .A3(new_n288), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n299), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n420), .A2(new_n423), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n328), .B(new_n354), .C1(new_n349), .C2(new_n346), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n469), .A2(new_n470), .A3(new_n336), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n469), .B2(new_n336), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n336), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n470), .A3(new_n336), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n317), .B2(new_n318), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n478), .A3(new_n362), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n367), .A2(new_n366), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n362), .B1(new_n482), .B2(new_n339), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n473), .A2(new_n478), .A3(KEYINPUT40), .A4(new_n362), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n465), .B1(new_n467), .B2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT85), .A3(new_n466), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT37), .B1(new_n401), .B2(new_n406), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n417), .A2(new_n492), .A3(new_n418), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n493), .A3(new_n410), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n411), .B1(new_n494), .B2(KEYINPUT38), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n364), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n483), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n371), .A2(new_n362), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT6), .B1(new_n357), .B2(new_n363), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n413), .A2(KEYINPUT38), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n403), .A2(new_n405), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n390), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n397), .A2(new_n400), .A3(new_n392), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n492), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n505), .B1(new_n504), .B2(new_n509), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n456), .B1(new_n502), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n464), .B1(new_n490), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n460), .A2(new_n455), .A3(new_n462), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT35), .B1(new_n515), .B2(new_n424), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n420), .A2(new_n517), .A3(new_n423), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(new_n501), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n462), .A2(new_n455), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n460), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(G29gat), .A2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n532));
  INV_X1    g331(.A(G36gat), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n532), .A2(KEYINPUT90), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT90), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n525), .A2(KEYINPUT89), .A3(KEYINPUT15), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n530), .A2(new_n536), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n532), .A2(new_n533), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n542), .A2(new_n531), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n524), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n541), .A2(KEYINPUT95), .A3(KEYINPUT17), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT92), .ZN(new_n551));
  INV_X1    g350(.A(G8gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n554));
  INV_X1    g353(.A(G1gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n552), .B1(new_n557), .B2(KEYINPUT94), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n553), .B(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n555), .A2(KEYINPUT16), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  OAI221_X1 g362(.A(new_n557), .B1(KEYINPUT94), .B2(new_n552), .C1(new_n560), .C2(new_n561), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n545), .A2(new_n566), .A3(new_n546), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n549), .A2(new_n551), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n545), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(KEYINPUT18), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n570), .B(new_n545), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n569), .B(KEYINPUT13), .Z(new_n579));
  AOI22_X1  g378(.A1(new_n576), .A2(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G169gat), .B(G197gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT12), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n574), .A2(new_n575), .A3(new_n580), .A4(new_n587), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n594));
  XOR2_X1   g393(.A(G57gat), .B(G64gat), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G71gat), .B(G78gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(new_n594), .A3(new_n596), .A4(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n565), .B1(new_n592), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n607), .B(new_n565), .C1(new_n592), .C2(new_n602), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT99), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n609), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n609), .B2(new_n610), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G99gat), .ZN(new_n620));
  INV_X1    g419(.A(G106gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  OAI21_X1  g425(.A(G92gat), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n627), .A2(new_n629), .B1(new_n625), .B2(new_n626), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT8), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n623), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n632), .B2(new_n623), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n624), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n634), .A3(new_n624), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n549), .A2(new_n551), .A3(new_n567), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n544), .B2(new_n541), .ZN(new_n642));
  NAND2_X1  g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT100), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(KEYINPUT41), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n641), .B1(new_n639), .B2(new_n646), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n650));
  XNOR2_X1  g449(.A(G134gat), .B(G162gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n646), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n640), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n652), .B1(new_n656), .B2(new_n647), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n619), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT102), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n653), .B1(new_n648), .B2(new_n649), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(new_n652), .A3(new_n647), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n619), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g466(.A(G230gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n431), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n637), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n602), .B1(new_n671), .B2(new_n635), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n636), .A2(new_n599), .A3(new_n601), .A4(new_n637), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(KEYINPUT103), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n638), .A2(new_n675), .A3(new_n602), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT10), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT10), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n670), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n674), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n669), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n667), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n680), .A2(new_n682), .A3(new_n667), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n684), .A2(KEYINPUT104), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT104), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n659), .A2(new_n664), .A3(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n523), .A2(new_n591), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n374), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT105), .B(G1gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1324gat));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  AND3_X1   g494(.A1(new_n690), .A2(new_n466), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT42), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n523), .A2(new_n591), .ZN(new_n699));
  INV_X1    g498(.A(new_n689), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G8gat), .B1(new_n701), .B2(new_n467), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT42), .ZN(new_n703));
  INV_X1    g502(.A(new_n696), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n697), .B1(new_n696), .B2(KEYINPUT42), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n698), .B1(new_n705), .B2(new_n706), .ZN(G1325gat));
  NAND2_X1  g506(.A1(new_n460), .A2(new_n462), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n701), .A2(G15gat), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n299), .A2(new_n463), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n299), .A2(KEYINPUT107), .A3(new_n463), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n701), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n715), .ZN(G1326gat));
  NAND2_X1  g515(.A1(new_n690), .A2(new_n456), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT108), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(new_n619), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n688), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n662), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n699), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(G29gat), .A3(new_n374), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(KEYINPUT45), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n512), .A2(new_n501), .A3(new_n495), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n488), .A2(KEYINPUT85), .A3(new_n466), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT85), .B1(new_n488), .B2(new_n466), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n455), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n457), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n299), .A2(KEYINPUT107), .A3(new_n463), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(new_n299), .B2(new_n463), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n516), .A2(new_n521), .A3(KEYINPUT110), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT110), .B1(new_n516), .B2(new_n521), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n734), .A2(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n662), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n514), .B2(new_n522), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n740), .A2(new_n744), .B1(new_n745), .B2(KEYINPUT44), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n591), .A2(new_n722), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n729), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n739), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n516), .A2(new_n521), .A3(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n714), .A2(new_n733), .A3(new_n457), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n743), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  INV_X1    g554(.A(new_n464), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n733), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n516), .A2(new_n521), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(new_n741), .ZN(new_n760));
  OAI211_X1 g559(.A(KEYINPUT112), .B(new_n747), .C1(new_n754), .C2(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n749), .A2(new_n691), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(G29gat), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n727), .B(new_n728), .C1(new_n762), .C2(new_n763), .ZN(G1328gat));
  NAND2_X1  g563(.A1(new_n466), .A2(new_n533), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT46), .B1(new_n725), .B2(new_n765), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n765), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n749), .A2(new_n466), .A3(new_n761), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n533), .ZN(G1329gat));
  NAND2_X1  g568(.A1(new_n740), .A2(new_n744), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n737), .A3(new_n747), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G43gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n725), .A2(G43gat), .A3(new_n708), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(KEYINPUT47), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n749), .A2(new_n737), .A3(new_n761), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(G43gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g579(.A1(new_n772), .A2(new_n456), .A3(new_n747), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G50gat), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n455), .A2(G50gat), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n782), .B(KEYINPUT48), .C1(new_n725), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n725), .A2(new_n783), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n749), .A2(new_n456), .A3(new_n761), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(G50gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g587(.A(new_n688), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n591), .A2(new_n659), .A3(new_n664), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n752), .B2(new_n753), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n691), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g592(.A(new_n467), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n799), .B(new_n801), .ZN(G1333gat));
  NAND2_X1  g601(.A1(new_n791), .A2(new_n737), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n708), .A2(G71gat), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n803), .A2(G71gat), .B1(new_n791), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n456), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g607(.A1(new_n589), .A2(new_n590), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n619), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n688), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n772), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G85gat), .B1(new_n813), .B2(new_n374), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n811), .A2(new_n662), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n740), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n789), .A2(new_n626), .A3(new_n691), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(G1336gat));
  XOR2_X1   g622(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n824));
  NAND3_X1  g623(.A1(new_n772), .A2(new_n466), .A3(new_n812), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(G92gat), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n467), .A2(G92gat), .A3(new_n688), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n818), .B2(new_n819), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n831), .B(new_n828), .C1(new_n818), .C2(new_n819), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n826), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n812), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n746), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n628), .B1(new_n835), .B2(new_n466), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT52), .B1(new_n836), .B2(new_n829), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(G1337gat));
  OAI21_X1  g637(.A(G99gat), .B1(new_n813), .B2(new_n714), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n789), .A2(new_n620), .A3(new_n460), .A4(new_n462), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n821), .B2(new_n840), .ZN(G1338gat));
  NAND3_X1  g640(.A1(new_n789), .A2(new_n456), .A3(new_n621), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT117), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n621), .B1(new_n835), .B2(new_n456), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT53), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G106gat), .B1(new_n813), .B2(new_n455), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n844), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(G1339gat));
  NOR2_X1   g650(.A1(new_n689), .A2(new_n809), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n677), .A2(new_n670), .A3(new_n679), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n680), .A3(KEYINPUT54), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(new_n670), .C1(new_n677), .C2(new_n679), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  INV_X1    g656(.A(new_n667), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT55), .B(new_n854), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n685), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n569), .B1(new_n568), .B2(new_n571), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n578), .A2(new_n579), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n586), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n862), .A2(new_n590), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n619), .B1(new_n869), .B2(new_n741), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n590), .B(new_n868), .C1(new_n686), .C2(new_n687), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n685), .A3(new_n861), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n662), .B(new_n871), .C1(new_n591), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n852), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n515), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n466), .A2(new_n374), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n591), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(G113gat), .Z(G1340gat));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n877), .A2(new_n688), .B1(new_n880), .B2(G120gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(G120gat), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(G1341gat));
  NOR2_X1   g682(.A1(new_n877), .A2(new_n721), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(new_n206), .ZN(G1342gat));
  NOR2_X1   g684(.A1(new_n874), .A2(new_n374), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n515), .A2(G134gat), .A3(new_n466), .A4(new_n662), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT120), .Z(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g690(.A(G134gat), .B1(new_n877), .B2(new_n662), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G1343gat));
  NOR3_X1   g692(.A1(new_n737), .A2(new_n874), .A3(new_n455), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n876), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n307), .A3(new_n809), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n714), .A2(KEYINPUT121), .A3(new_n876), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT121), .B1(new_n714), .B2(new_n876), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n871), .A2(new_n662), .ZN(new_n900));
  INV_X1    g699(.A(new_n872), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n809), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n590), .A2(new_n868), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n741), .B1(new_n872), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n721), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n902), .A2(new_n905), .B1(new_n809), .B2(new_n689), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(KEYINPUT57), .A3(new_n456), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n874), .B2(new_n455), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n899), .A2(new_n809), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n896), .B1(new_n912), .B2(new_n307), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT58), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n896), .C1(new_n912), .C2(new_n307), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1344gat));
  NAND3_X1  g716(.A1(new_n895), .A2(new_n309), .A3(new_n789), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n910), .B(new_n789), .C1(new_n898), .C2(new_n897), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(G148gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(G148gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT122), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n918), .B(new_n925), .C1(new_n921), .C2(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(G155gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n895), .A2(new_n928), .A3(new_n619), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n899), .A2(new_n619), .A3(new_n910), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n929), .B1(new_n931), .B2(new_n928), .ZN(G1346gat));
  NOR4_X1   g731(.A1(new_n466), .A2(new_n455), .A3(G162gat), .A4(new_n662), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n886), .A2(new_n714), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n899), .A2(new_n741), .A3(new_n910), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(G162gat), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(G1347gat));
  OAI21_X1  g737(.A(KEYINPUT124), .B1(new_n515), .B2(new_n467), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n515), .A2(KEYINPUT124), .A3(new_n467), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(new_n691), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n906), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n809), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n467), .A2(new_n691), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n874), .A2(new_n515), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n809), .A2(G169gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1348gat));
  INV_X1    g747(.A(new_n946), .ZN(new_n949));
  OAI21_X1  g748(.A(G176gat), .B1(new_n949), .B2(new_n688), .ZN(new_n950));
  INV_X1    g749(.A(G176gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n942), .A2(new_n951), .A3(new_n789), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1349gat));
  NAND3_X1  g752(.A1(new_n942), .A2(new_n216), .A3(new_n619), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT125), .Z(new_n955));
  OAI21_X1  g754(.A(G183gat), .B1(new_n949), .B2(new_n721), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n959), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n949), .B2(new_n662), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n965), .B1(KEYINPUT126), .B2(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n964), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n942), .A2(new_n215), .A3(new_n741), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G1351gat));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n737), .A2(new_n945), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n910), .A2(new_n809), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n972), .B2(KEYINPUT127), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n973), .B1(KEYINPUT127), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n894), .A2(new_n944), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n970), .A3(new_n809), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n974), .A2(new_n977), .ZN(G1352gat));
  OR3_X1    g777(.A1(new_n975), .A2(G204gat), .A3(new_n688), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n910), .A2(new_n971), .ZN(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n981), .B2(new_n688), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(G1353gat));
  OR3_X1    g783(.A1(new_n975), .A2(G211gat), .A3(new_n721), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n910), .A2(new_n619), .A3(new_n971), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  OR3_X1    g788(.A1(new_n975), .A2(G218gat), .A3(new_n662), .ZN(new_n990));
  OAI21_X1  g789(.A(G218gat), .B1(new_n981), .B2(new_n662), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


