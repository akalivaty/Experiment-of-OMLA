//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1118;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n461), .A2(new_n463), .B1(new_n464), .B2(G101), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(G160));
  XNOR2_X1  g043(.A(new_n461), .B(KEYINPUT68), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(new_n462), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G124), .ZN(new_n471));
  OR2_X1    g046(.A1(G100), .A2(G2105), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n472), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(G136), .B2(new_n475), .ZN(G162));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(G114), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g055(.A1(G102), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n461), .B2(new_n488), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n485), .B(new_n486), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n491), .A2(new_n490), .ZN(new_n498));
  NAND2_X1  g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n488), .B1(new_n491), .B2(new_n490), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n502), .B2(new_n492), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(new_n485), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n497), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n510), .B2(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(G651), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n510), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n507), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(G88), .B1(new_n523), .B2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  XNOR2_X1  g101(.A(new_n523), .B(KEYINPUT73), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n519), .A2(new_n520), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G89), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(G63), .B2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n528), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(new_n522), .A2(G90), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n527), .B2(G52), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n518), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n543), .A2(G651), .B1(new_n522), .B2(G81), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n523), .B(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g126(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(G188));
  NAND3_X1  g131(.A1(new_n531), .A2(G53), .A3(G543), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n522), .A2(G91), .ZN(new_n560));
  INV_X1    g135(.A(new_n509), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT5), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G65), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n560), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n559), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n522), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n523), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n508), .B2(new_n509), .ZN(new_n578));
  AND2_X1   g153(.A1(G73), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n531), .A2(G86), .A3(new_n510), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n531), .A2(G48), .A3(G543), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G305));
  XNOR2_X1  g158(.A(KEYINPUT78), .B(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n527), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n518), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n522), .B2(G85), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n522), .A2(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n518), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n527), .A2(G54), .B1(G651), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n549), .ZN(G323));
  XOR2_X1   g188(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n614));
  XNOR2_X1  g189(.A(G323), .B(new_n614), .ZN(G282));
  NAND2_X1  g190(.A1(new_n461), .A2(new_n464), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n475), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n470), .A2(G123), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(G2096), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n626), .A3(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2430), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT82), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n630), .B2(new_n631), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(new_n643), .A3(G14), .ZN(G401));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n658), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n658), .B2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n672), .B(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G6), .A2(G16), .ZN(new_n679));
  INV_X1    g254(.A(G305), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(G16), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT32), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1981), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT89), .Z(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n684), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(G1971), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(G1971), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n684), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  NOR4_X1   g269(.A1(new_n683), .A2(new_n688), .A3(new_n689), .A4(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  OR2_X1    g273(.A1(G25), .A2(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n475), .A2(G131), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n462), .A2(G107), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n470), .A2(KEYINPUT87), .A3(G119), .ZN(new_n703));
  AOI21_X1  g278(.A(KEYINPUT87), .B1(new_n470), .B2(G119), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n700), .B1(new_n701), .B2(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n699), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT35), .B(G1991), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT88), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(G16), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  INV_X1    g288(.A(new_n710), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n697), .A2(new_n698), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT36), .Z(new_n717));
  NOR2_X1   g292(.A1(G168), .A2(new_n684), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n684), .B2(G21), .ZN(new_n719));
  INV_X1    g294(.A(G1966), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  NAND2_X1  g296(.A1(G171), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G5), .B2(G16), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n721), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n724), .B(new_n725), .C1(new_n720), .C2(new_n719), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n706), .A2(G33), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n462), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G139), .B2(new_n475), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n706), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT93), .Z(new_n735));
  AOI21_X1  g310(.A(new_n726), .B1(G2072), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G35), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G162), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT29), .B(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G19), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n549), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1341), .ZN(new_n743));
  INV_X1    g318(.A(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n745), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n625), .B2(new_n706), .ZN(new_n750));
  INV_X1    g325(.A(G34), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT24), .B2(new_n751), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n467), .B2(new_n706), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n740), .A2(new_n743), .A3(new_n750), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n684), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT23), .ZN(new_n759));
  INV_X1    g334(.A(G299), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n684), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1956), .Z(new_n762));
  NOR2_X1   g337(.A1(G4), .A2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT90), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n601), .B2(new_n684), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1348), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n736), .A2(new_n757), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n706), .A2(G32), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n475), .A2(G141), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n470), .A2(G129), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G105), .B2(new_n464), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(new_n706), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n735), .A2(G2072), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n706), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n706), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G2078), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n706), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n475), .A2(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n470), .A2(G128), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n462), .A2(G116), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n780), .A2(new_n781), .A3(new_n784), .A4(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n717), .A2(new_n767), .A3(new_n795), .ZN(G311));
  INV_X1    g371(.A(G311), .ZN(G150));
  NAND2_X1  g372(.A1(new_n602), .A2(G559), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT38), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n548), .B(KEYINPUT97), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n537), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G55), .B2(new_n527), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n522), .A2(G93), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n800), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n799), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  AOI21_X1  g389(.A(G860), .B1(new_n812), .B2(KEYINPUT39), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n808), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(G145));
  XNOR2_X1  g394(.A(new_n792), .B(new_n775), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(new_n495), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n495), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n733), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n733), .A2(new_n823), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n705), .B(new_n617), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(G118), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(KEYINPUT101), .B1(new_n829), .B2(G2105), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT101), .B2(new_n828), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n470), .A2(G130), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n475), .A2(new_n833), .A3(G142), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n475), .B2(G142), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n831), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n827), .B(new_n836), .Z(new_n837));
  OR2_X1    g412(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n826), .A2(new_n837), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n625), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G162), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n840), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g420(.A1(new_n808), .A2(new_n605), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n811), .B(new_n611), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n601), .B(new_n760), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT41), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n853), .B2(new_n847), .ZN(new_n854));
  XNOR2_X1  g429(.A(G290), .B(G305), .ZN(new_n855));
  XNOR2_X1  g430(.A(G303), .B(G288), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n855), .B(new_n856), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT42), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n854), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n846), .B1(new_n860), .B2(new_n605), .ZN(G295));
  OAI21_X1  g436(.A(new_n846), .B1(new_n860), .B2(new_n605), .ZN(G331));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  XNOR2_X1  g438(.A(G168), .B(G171), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n811), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n809), .A2(new_n810), .A3(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n848), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n851), .A2(new_n852), .B1(new_n867), .B2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n857), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n869), .B(new_n857), .C1(new_n870), .C2(new_n871), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT43), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n879), .B(new_n857), .C1(new_n870), .C2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n874), .A2(new_n881), .A3(new_n882), .A4(new_n875), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n863), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI211_X1 g461(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n878), .C2(new_n883), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n877), .A2(KEYINPUT43), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n874), .A2(new_n881), .A3(new_n875), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT44), .B1(new_n889), .B2(new_n882), .ZN(new_n890));
  OAI22_X1  g465(.A1(new_n886), .A2(new_n887), .B1(new_n888), .B2(new_n890), .ZN(G397));
  INV_X1    g466(.A(G1384), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n497), .B2(new_n504), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT50), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n495), .A2(new_n892), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(KEYINPUT50), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n495), .A2(new_n496), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n503), .A2(KEYINPUT70), .A3(new_n485), .ZN(new_n899));
  AOI21_X1  g474(.A(G1384), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT50), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G40), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n467), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n895), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT115), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT115), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n895), .A2(new_n902), .A3(new_n907), .A4(new_n904), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT121), .B(G1961), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g486(.A1(G160), .A2(G40), .ZN(new_n912));
  AOI21_X1  g487(.A(G1384), .B1(new_n503), .B2(new_n485), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(KEYINPUT45), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(KEYINPUT45), .B2(new_n900), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n911), .B1(new_n915), .B2(G2078), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n912), .B1(new_n917), .B2(new_n896), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT122), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT53), .B1(new_n919), .B2(G2078), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n919), .B2(G2078), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n918), .B(new_n921), .C1(new_n917), .C2(new_n896), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n910), .A2(new_n916), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G171), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n893), .B2(new_n917), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n925), .A2(new_n911), .A3(G2078), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n910), .A2(G301), .A3(new_n916), .A4(new_n926), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT123), .A2(new_n924), .A3(KEYINPUT54), .A4(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT54), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n923), .B2(G171), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT123), .B1(new_n930), .B2(new_n927), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n912), .A2(new_n896), .ZN(new_n933));
  INV_X1    g508(.A(G8), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n573), .A2(new_n575), .A3(G1976), .A4(new_n574), .ZN(new_n936));
  INV_X1    g511(.A(G1976), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT52), .B1(G288), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n581), .A2(new_n582), .ZN(new_n940));
  INV_X1    g515(.A(G1981), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n940), .B(new_n580), .C1(KEYINPUT108), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n580), .B2(KEYINPUT108), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G305), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT49), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(KEYINPUT49), .A3(new_n944), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n935), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(G8), .B(new_n936), .C1(new_n912), .C2(new_n896), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n950), .A2(KEYINPUT107), .A3(KEYINPUT52), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT107), .B1(new_n950), .B2(KEYINPUT52), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n939), .B(new_n949), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n912), .B1(KEYINPUT50), .B2(new_n896), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n901), .B(new_n892), .C1(new_n497), .C2(new_n504), .ZN(new_n955));
  INV_X1    g530(.A(G2090), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n904), .B1(new_n896), .B2(new_n917), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n893), .B2(new_n917), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n959), .B2(G1971), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G8), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(G8), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT55), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n953), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n895), .A2(new_n902), .A3(new_n956), .A4(new_n904), .ZN(new_n965));
  INV_X1    g540(.A(G1971), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n915), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n934), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n963), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n895), .A2(new_n902), .A3(new_n755), .A4(new_n904), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n925), .A2(new_n720), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n934), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n975));
  NOR2_X1   g550(.A1(G168), .A2(new_n934), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(KEYINPUT51), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n976), .B(KEYINPUT119), .Z(new_n979));
  OAI21_X1  g554(.A(KEYINPUT51), .B1(new_n979), .B2(new_n974), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n974), .B2(new_n977), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n973), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n976), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n971), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n910), .A2(new_n916), .A3(new_n926), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n986), .A2(G171), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n923), .A2(G171), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n929), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n932), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1348), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n906), .A2(new_n992), .A3(new_n908), .ZN(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n933), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT116), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n760), .A2(KEYINPUT57), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n569), .A2(KEYINPUT113), .ZN(new_n1001));
  INV_X1    g576(.A(new_n559), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n560), .B(new_n1003), .C1(new_n567), .C2(new_n568), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT114), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1005), .A2(KEYINPUT114), .A3(new_n1007), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT56), .B(G2072), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n914), .B(new_n1012), .C1(KEYINPUT45), .C2(new_n900), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n954), .A2(new_n955), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(G1956), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(new_n601), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n997), .A2(new_n999), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1013), .B(KEYINPUT117), .C1(new_n1014), .C2(G1956), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1011), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n993), .A2(new_n998), .A3(new_n995), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n998), .B1(new_n993), .B2(new_n995), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT60), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT60), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n997), .A2(new_n1028), .A3(new_n999), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1027), .A2(new_n1029), .A3(new_n602), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT61), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n760), .A2(KEYINPUT57), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1010), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n1008), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1956), .B1(new_n954), .B2(new_n955), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n959), .B2(new_n1012), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1031), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1022), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT58), .B(G1341), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n915), .A2(G1996), .B1(new_n933), .B2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1040), .A2(KEYINPUT59), .A3(new_n549), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT59), .B1(new_n1040), .B2(new_n549), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n1045));
  NOR2_X1   g620(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1016), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1044), .B(new_n1047), .C1(new_n1027), .C2(new_n602), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1024), .B1(new_n1030), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n991), .A2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n934), .B(G286), .C1(new_n972), .C2(new_n973), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n964), .A2(new_n970), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n964), .A2(KEYINPUT110), .A3(new_n970), .A4(new_n1051), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT111), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1056), .A4(new_n1055), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1056), .B(new_n953), .C1(new_n969), .C2(new_n968), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(new_n1051), .C1(new_n969), .C2(new_n968), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n970), .A2(new_n953), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n935), .B(KEYINPUT109), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n949), .A2(new_n937), .A3(new_n691), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n680), .A2(new_n941), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1050), .A2(KEYINPUT124), .A3(new_n1064), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1047), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1028), .B1(new_n997), .B2(new_n999), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n601), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1027), .A2(new_n1029), .A3(new_n602), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1023), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n989), .B(new_n985), .C1(new_n928), .C2(new_n931), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1064), .B(new_n1070), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n982), .A2(new_n984), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1082));
  INV_X1    g657(.A(new_n987), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1082), .A2(new_n971), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(KEYINPUT62), .B2(new_n1081), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1071), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n896), .A2(new_n917), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(new_n912), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n705), .A2(new_n710), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n792), .B(new_n994), .ZN(new_n1090));
  INV_X1    g665(.A(G1996), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n775), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n705), .A2(new_n710), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(G290), .B(G1986), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1088), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1086), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1088), .ZN(new_n1098));
  NOR4_X1   g673(.A1(G290), .A2(new_n1087), .A3(G1986), .A4(new_n912), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT48), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1101));
  OAI22_X1  g676(.A1(new_n1101), .A2(new_n1089), .B1(G2067), .B2(new_n792), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1098), .A2(new_n1100), .B1(new_n1102), .B2(new_n1088), .ZN(new_n1103));
  NAND2_X1  g678(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1104));
  NOR4_X1   g679(.A1(new_n1087), .A2(new_n912), .A3(G1996), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1090), .A2(new_n776), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1088), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT126), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1088), .B(new_n1091), .C1(KEYINPUT125), .C2(KEYINPUT46), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1105), .B(new_n1108), .C1(new_n1104), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT47), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1103), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1113), .B2(new_n1112), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1097), .A2(new_n1115), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g691(.A1(G401), .A2(new_n459), .A3(G227), .A4(G229), .ZN(new_n1118));
  NAND3_X1  g692(.A1(new_n844), .A2(new_n884), .A3(new_n1118), .ZN(G225));
  INV_X1    g693(.A(G225), .ZN(G308));
endmodule


