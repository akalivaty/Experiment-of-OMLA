

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n907), .A2(n687), .ZN(n693) );
  NOR2_X1 U553 ( .A1(G299), .A2(n703), .ZN(n700) );
  NOR2_X1 U554 ( .A1(n920), .A2(n686), .ZN(n687) );
  XNOR2_X2 U555 ( .A(n537), .B(KEYINPUT65), .ZN(n605) );
  XNOR2_X1 U556 ( .A(n708), .B(n707), .ZN(n714) );
  AND2_X1 U557 ( .A1(n749), .A2(n746), .ZN(n747) );
  XOR2_X1 U558 ( .A(KEYINPUT14), .B(n555), .Z(n519) );
  INV_X1 U559 ( .A(KEYINPUT27), .ZN(n694) );
  XNOR2_X1 U560 ( .A(n695), .B(n694), .ZN(n698) );
  INV_X1 U561 ( .A(KEYINPUT90), .ZN(n699) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n707) );
  NOR2_X1 U563 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U564 ( .A(n681), .B(n680), .ZN(n710) );
  INV_X1 U565 ( .A(n936), .ZN(n745) );
  NOR2_X1 U566 ( .A1(n745), .A2(KEYINPUT33), .ZN(n746) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n756) );
  NAND2_X1 U568 ( .A1(n748), .A2(n747), .ZN(n753) );
  INV_X1 U569 ( .A(G651), .ZN(n524) );
  NAND2_X1 U570 ( .A1(n888), .A2(G138), .ZN(n558) );
  INV_X1 U571 ( .A(KEYINPUT17), .ZN(n532) );
  AND2_X2 U572 ( .A1(n538), .A2(G2104), .ZN(n887) );
  OR2_X1 U573 ( .A1(n801), .A2(n800), .ZN(n819) );
  NOR2_X1 U574 ( .A1(G651), .A2(n624), .ZN(n647) );
  AND2_X1 U575 ( .A1(n564), .A2(n563), .ZN(G164) );
  XOR2_X1 U576 ( .A(KEYINPUT70), .B(n557), .Z(n920) );
  NOR2_X1 U577 ( .A1(n542), .A2(n541), .ZN(G160) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U579 ( .A1(n639), .A2(G91), .ZN(n520) );
  XOR2_X1 U580 ( .A(KEYINPUT67), .B(n520), .Z(n522) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n624) );
  NOR2_X1 U582 ( .A1(n624), .A2(n524), .ZN(n640) );
  NAND2_X1 U583 ( .A1(n640), .A2(G78), .ZN(n521) );
  NAND2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U585 ( .A(KEYINPUT68), .B(n523), .ZN(n529) );
  NOR2_X1 U586 ( .A1(G543), .A2(n524), .ZN(n525) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n525), .Z(n526) );
  XNOR2_X2 U588 ( .A(KEYINPUT66), .B(n526), .ZN(n643) );
  NAND2_X1 U589 ( .A1(G65), .A2(n643), .ZN(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT69), .B(n527), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n647), .A2(G53), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(G299) );
  NOR2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XNOR2_X2 U595 ( .A(n533), .B(n532), .ZN(n888) );
  NAND2_X1 U596 ( .A1(n888), .A2(G137), .ZN(n536) );
  INV_X1 U597 ( .A(G2105), .ZN(n538) );
  NAND2_X1 U598 ( .A1(G101), .A2(n887), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(n534), .Z(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  NAND2_X1 U602 ( .A1(G113), .A2(n605), .ZN(n540) );
  NOR2_X2 U603 ( .A1(G2104), .A2(n538), .ZN(n892) );
  NAND2_X1 U604 ( .A1(G125), .A2(n892), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U606 ( .A1(G85), .A2(n639), .ZN(n544) );
  NAND2_X1 U607 ( .A1(G72), .A2(n640), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G47), .A2(n647), .ZN(n546) );
  NAND2_X1 U610 ( .A1(G60), .A2(n643), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(G290) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G860), .ZN(n599) );
  NAND2_X1 U615 ( .A1(n639), .A2(G81), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT12), .ZN(n551) );
  NAND2_X1 U617 ( .A1(G68), .A2(n640), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT13), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G43), .A2(n647), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n643), .A2(G56), .ZN(n555) );
  NOR2_X1 U623 ( .A1(n556), .A2(n519), .ZN(n557) );
  OR2_X1 U624 ( .A1(n599), .A2(n920), .ZN(G153) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U628 ( .A(n558), .B(KEYINPUT84), .ZN(n564) );
  AND2_X1 U629 ( .A1(n887), .A2(G102), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G114), .A2(n605), .ZN(n560) );
  NAND2_X1 U631 ( .A1(G126), .A2(n892), .ZN(n559) );
  NAND2_X1 U632 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U634 ( .A1(G52), .A2(n647), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G64), .A2(n643), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G90), .A2(n639), .ZN(n568) );
  NAND2_X1 U638 ( .A1(G77), .A2(n640), .ZN(n567) );
  NAND2_X1 U639 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U641 ( .A1(n571), .A2(n570), .ZN(G171) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n822) );
  NAND2_X1 U645 ( .A1(n822), .A2(G567), .ZN(n573) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n640), .A2(G79), .ZN(n574) );
  XOR2_X1 U650 ( .A(KEYINPUT71), .B(n574), .Z(n576) );
  NAND2_X1 U651 ( .A1(n647), .A2(G54), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U653 ( .A(KEYINPUT72), .B(n577), .ZN(n581) );
  NAND2_X1 U654 ( .A1(G92), .A2(n639), .ZN(n579) );
  NAND2_X1 U655 ( .A1(G66), .A2(n643), .ZN(n578) );
  NAND2_X1 U656 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n582), .Z(n907) );
  INV_X1 U659 ( .A(n907), .ZN(n922) );
  INV_X1 U660 ( .A(G868), .ZN(n650) );
  NAND2_X1 U661 ( .A1(n922), .A2(n650), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(G284) );
  XNOR2_X1 U663 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G51), .A2(n647), .ZN(n586) );
  NAND2_X1 U665 ( .A1(G63), .A2(n643), .ZN(n585) );
  NAND2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U667 ( .A(n588), .B(n587), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n639), .A2(G89), .ZN(n589) );
  XNOR2_X1 U669 ( .A(n589), .B(KEYINPUT4), .ZN(n591) );
  NAND2_X1 U670 ( .A1(G76), .A2(n640), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U672 ( .A(KEYINPUT5), .B(n592), .ZN(n593) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(n593), .ZN(n594) );
  NOR2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U675 ( .A(KEYINPUT7), .B(n596), .Z(G168) );
  XOR2_X1 U676 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U677 ( .A1(G286), .A2(n650), .ZN(n598) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U679 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n600), .A2(n907), .ZN(n601) );
  XNOR2_X1 U682 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(n920), .A2(G868), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n907), .A2(G868), .ZN(n602) );
  NOR2_X1 U685 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G111), .A2(n605), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G99), .A2(n887), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G135), .A2(n888), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n892), .A2(G123), .ZN(n608) );
  XOR2_X1 U692 ( .A(KEYINPUT18), .B(n608), .Z(n609) );
  NOR2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT75), .ZN(n1005) );
  XNOR2_X1 U696 ( .A(n1005), .B(G2096), .ZN(n615) );
  INV_X1 U697 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G559), .A2(n907), .ZN(n616) );
  XNOR2_X1 U700 ( .A(n616), .B(n920), .ZN(n659) );
  NOR2_X1 U701 ( .A1(G860), .A2(n659), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G93), .A2(n639), .ZN(n618) );
  NAND2_X1 U703 ( .A1(G80), .A2(n640), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U705 ( .A1(G55), .A2(n647), .ZN(n620) );
  NAND2_X1 U706 ( .A1(G67), .A2(n643), .ZN(n619) );
  NAND2_X1 U707 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n652) );
  XOR2_X1 U709 ( .A(n623), .B(n652), .Z(G145) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G49), .A2(n647), .ZN(n626) );
  NAND2_X1 U712 ( .A1(G87), .A2(n624), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U714 ( .A1(n643), .A2(n627), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U716 ( .A(n630), .B(KEYINPUT76), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G86), .A2(n639), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G48), .A2(n647), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G73), .A2(n640), .ZN(n633) );
  XNOR2_X1 U721 ( .A(n633), .B(KEYINPUT77), .ZN(n634) );
  XNOR2_X1 U722 ( .A(n634), .B(KEYINPUT2), .ZN(n635) );
  NOR2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U724 ( .A1(G61), .A2(n643), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G88), .A2(n639), .ZN(n642) );
  NAND2_X1 U727 ( .A1(G75), .A2(n640), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n643), .A2(G62), .ZN(n644) );
  XOR2_X1 U730 ( .A(KEYINPUT78), .B(n644), .Z(n645) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n647), .A2(G50), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  NAND2_X1 U735 ( .A1(n650), .A2(n652), .ZN(n651) );
  XNOR2_X1 U736 ( .A(n651), .B(KEYINPUT80), .ZN(n662) );
  XOR2_X1 U737 ( .A(n652), .B(G305), .Z(n655) );
  XNOR2_X1 U738 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U739 ( .A(n653), .B(G290), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U741 ( .A(G288), .B(n656), .ZN(n658) );
  XNOR2_X1 U742 ( .A(G299), .B(G166), .ZN(n657) );
  XNOR2_X1 U743 ( .A(n658), .B(n657), .ZN(n904) );
  XNOR2_X1 U744 ( .A(n904), .B(n659), .ZN(n660) );
  NAND2_X1 U745 ( .A1(G868), .A2(n660), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U747 ( .A(KEYINPUT81), .B(n663), .Z(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n664) );
  XNOR2_X1 U750 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n669) );
  XNOR2_X1 U756 ( .A(KEYINPUT22), .B(n669), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n670), .A2(G96), .ZN(n671) );
  NOR2_X1 U758 ( .A1(n671), .A2(G218), .ZN(n672) );
  XNOR2_X1 U759 ( .A(n672), .B(KEYINPUT83), .ZN(n828) );
  NAND2_X1 U760 ( .A1(n828), .A2(G2106), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n673) );
  NOR2_X1 U762 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U763 ( .A1(G108), .A2(n674), .ZN(n827) );
  NAND2_X1 U764 ( .A1(n827), .A2(G567), .ZN(n675) );
  NAND2_X1 U765 ( .A1(n676), .A2(n675), .ZN(n916) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U767 ( .A1(n916), .A2(n677), .ZN(n826) );
  NAND2_X1 U768 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n755) );
  INV_X1 U770 ( .A(n755), .ZN(n679) );
  NAND2_X1 U771 ( .A1(n679), .A2(n756), .ZN(n681) );
  INV_X1 U772 ( .A(KEYINPUT64), .ZN(n680) );
  INV_X1 U773 ( .A(n710), .ZN(n717) );
  INV_X1 U774 ( .A(G1996), .ZN(n972) );
  NOR2_X1 U775 ( .A1(n717), .A2(n972), .ZN(n683) );
  XNOR2_X1 U776 ( .A(KEYINPUT26), .B(KEYINPUT89), .ZN(n682) );
  XNOR2_X1 U777 ( .A(n683), .B(n682), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n717), .A2(G1341), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U780 ( .A1(n907), .A2(n687), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n710), .B(KEYINPUT88), .ZN(n696) );
  NAND2_X1 U782 ( .A1(n696), .A2(G2067), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n717), .A2(G1348), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n702) );
  NAND2_X1 U787 ( .A1(n696), .A2(G2072), .ZN(n695) );
  INV_X1 U788 ( .A(n696), .ZN(n709) );
  NAND2_X1 U789 ( .A1(G1956), .A2(n709), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n703) );
  XNOR2_X1 U791 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U793 ( .A1(G299), .A2(n703), .ZN(n704) );
  XNOR2_X1 U794 ( .A(n704), .B(KEYINPUT28), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n708) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .Z(n973) );
  NOR2_X1 U797 ( .A1(n973), .A2(n709), .ZN(n712) );
  NOR2_X1 U798 ( .A1(G1961), .A2(n710), .ZN(n711) );
  NOR2_X1 U799 ( .A1(n712), .A2(n711), .ZN(n715) );
  OR2_X1 U800 ( .A1(n715), .A2(G301), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n725) );
  NAND2_X1 U802 ( .A1(n715), .A2(G301), .ZN(n716) );
  XNOR2_X1 U803 ( .A(n716), .B(KEYINPUT91), .ZN(n722) );
  NAND2_X1 U804 ( .A1(n717), .A2(G8), .ZN(n809) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n809), .ZN(n738) );
  NOR2_X1 U806 ( .A1(n717), .A2(G2084), .ZN(n735) );
  NOR2_X1 U807 ( .A1(n738), .A2(n735), .ZN(n718) );
  NAND2_X1 U808 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n720), .A2(G168), .ZN(n721) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n723), .Z(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n736) );
  NAND2_X1 U813 ( .A1(n736), .A2(G286), .ZN(n726) );
  XNOR2_X1 U814 ( .A(n726), .B(KEYINPUT92), .ZN(n732) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n809), .ZN(n728) );
  NOR2_X1 U816 ( .A1(n717), .A2(G2090), .ZN(n727) );
  NOR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n729), .A2(G303), .ZN(n730) );
  XOR2_X1 U819 ( .A(KEYINPUT93), .B(n730), .Z(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n733), .A2(G8), .ZN(n734) );
  XNOR2_X1 U822 ( .A(n734), .B(KEYINPUT32), .ZN(n742) );
  NAND2_X1 U823 ( .A1(G8), .A2(n735), .ZN(n740) );
  INV_X1 U824 ( .A(n736), .ZN(n737) );
  NOR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n804) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n750), .A2(n743), .ZN(n933) );
  NAND2_X1 U831 ( .A1(n804), .A2(n933), .ZN(n744) );
  XNOR2_X1 U832 ( .A(n744), .B(KEYINPUT94), .ZN(n748) );
  INV_X1 U833 ( .A(n809), .ZN(n749) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n936) );
  NAND2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U838 ( .A(n754), .B(KEYINPUT95), .ZN(n801) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n917) );
  NOR2_X1 U840 ( .A1(n756), .A2(n755), .ZN(n796) );
  NAND2_X1 U841 ( .A1(n887), .A2(G104), .ZN(n757) );
  XOR2_X1 U842 ( .A(KEYINPUT85), .B(n757), .Z(n759) );
  NAND2_X1 U843 ( .A1(n888), .A2(G140), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U845 ( .A(KEYINPUT34), .B(n760), .ZN(n766) );
  NAND2_X1 U846 ( .A1(n892), .A2(G128), .ZN(n761) );
  XNOR2_X1 U847 ( .A(n761), .B(KEYINPUT86), .ZN(n763) );
  NAND2_X1 U848 ( .A1(G116), .A2(n605), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U850 ( .A(KEYINPUT35), .B(n764), .Z(n765) );
  NOR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U852 ( .A(KEYINPUT36), .B(n767), .ZN(n901) );
  XNOR2_X1 U853 ( .A(G2067), .B(KEYINPUT37), .ZN(n768) );
  NOR2_X1 U854 ( .A1(n901), .A2(n768), .ZN(n1002) );
  NAND2_X1 U855 ( .A1(n796), .A2(n1002), .ZN(n813) );
  AND2_X1 U856 ( .A1(n917), .A2(n813), .ZN(n799) );
  NAND2_X1 U857 ( .A1(n901), .A2(n768), .ZN(n769) );
  XNOR2_X1 U858 ( .A(KEYINPUT98), .B(n769), .ZN(n1014) );
  NAND2_X1 U859 ( .A1(n887), .A2(G105), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT38), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G141), .A2(n888), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G117), .A2(n605), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G129), .A2(n892), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n881) );
  AND2_X1 U867 ( .A1(n972), .A2(n881), .ZN(n997) );
  NAND2_X1 U868 ( .A1(G95), .A2(n887), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G131), .A2(n888), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G107), .A2(n605), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G119), .A2(n892), .ZN(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n882) );
  INV_X1 U875 ( .A(G1991), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n882), .A2(n785), .ZN(n784) );
  NOR2_X1 U877 ( .A1(n972), .A2(n881), .ZN(n783) );
  NOR2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n795) );
  INV_X1 U879 ( .A(n795), .ZN(n1000) );
  NOR2_X1 U880 ( .A1(G1986), .A2(G290), .ZN(n787) );
  AND2_X1 U881 ( .A1(n785), .A2(n882), .ZN(n786) );
  XNOR2_X1 U882 ( .A(KEYINPUT96), .B(n786), .ZN(n1001) );
  NOR2_X1 U883 ( .A1(n787), .A2(n1001), .ZN(n788) );
  XOR2_X1 U884 ( .A(KEYINPUT97), .B(n788), .Z(n789) );
  NOR2_X1 U885 ( .A1(n1000), .A2(n789), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n997), .A2(n790), .ZN(n791) );
  XNOR2_X1 U887 ( .A(n791), .B(KEYINPUT39), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n792), .A2(n813), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n1014), .A2(n793), .ZN(n794) );
  AND2_X1 U890 ( .A1(n794), .A2(n796), .ZN(n814) );
  XOR2_X1 U891 ( .A(G1986), .B(G290), .Z(n931) );
  NAND2_X1 U892 ( .A1(n795), .A2(n931), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U894 ( .A1(n814), .A2(n798), .ZN(n817) );
  NAND2_X1 U895 ( .A1(n799), .A2(n817), .ZN(n800) );
  NOR2_X1 U896 ( .A1(G2090), .A2(G303), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G8), .A2(n802), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n805), .A2(n809), .ZN(n811) );
  NOR2_X1 U900 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n806), .B(KEYINPUT24), .ZN(n807) );
  XNOR2_X1 U902 ( .A(KEYINPUT87), .B(n807), .ZN(n808) );
  OR2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n815) );
  OR2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n819), .A2(n818), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n820) );
  XNOR2_X1 U910 ( .A(n821), .B(n820), .ZN(G329) );
  NAND2_X1 U911 ( .A1(n822), .A2(G2106), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT103), .B(n823), .Z(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT104), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U924 ( .A(G2427), .B(G2443), .ZN(n839) );
  XOR2_X1 U925 ( .A(G2430), .B(KEYINPUT101), .Z(n831) );
  XNOR2_X1 U926 ( .A(G2454), .B(G2435), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U928 ( .A(G2438), .B(KEYINPUT100), .Z(n833) );
  XNOR2_X1 U929 ( .A(G1341), .B(G1348), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U931 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2446), .B(G2451), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n840), .A2(G14), .ZN(n841) );
  XOR2_X1 U936 ( .A(KEYINPUT102), .B(n841), .Z(G401) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n843) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT105), .B(G1991), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1981), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U949 ( .A(n852), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U950 ( .A(G1976), .B(G1986), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U952 ( .A(G1971), .B(G1956), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1961), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT106), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G136), .A2(n888), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n861), .B(KEYINPUT108), .ZN(n865) );
  XOR2_X1 U960 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n863) );
  NAND2_X1 U961 ( .A1(G124), .A2(n892), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G100), .A2(n887), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G112), .A2(n605), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G118), .A2(n605), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G130), .A2(n892), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G106), .A2(n887), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G142), .A2(n888), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT109), .B(n874), .ZN(n875) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n875), .ZN(n876) );
  NOR2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U977 ( .A(n878), .B(G162), .Z(n880) );
  XNOR2_X1 U978 ( .A(G164), .B(n1005), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(n886) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(n886), .B(n885), .Z(n900) );
  NAND2_X1 U984 ( .A1(G103), .A2(n887), .ZN(n890) );
  NAND2_X1 U985 ( .A1(G139), .A2(n888), .ZN(n889) );
  NAND2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U987 ( .A1(n605), .A2(G115), .ZN(n891) );
  XNOR2_X1 U988 ( .A(KEYINPUT111), .B(n891), .ZN(n895) );
  NAND2_X1 U989 ( .A1(n892), .A2(G127), .ZN(n893) );
  XOR2_X1 U990 ( .A(KEYINPUT110), .B(n893), .Z(n894) );
  NOR2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n896), .B(KEYINPUT47), .ZN(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n1010) );
  XNOR2_X1 U994 ( .A(G160), .B(n1010), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U996 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(n904), .Z(n906) );
  XNOR2_X1 U999 ( .A(G171), .B(n920), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(G286), .B(n907), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n910), .ZN(G397) );
  OR2_X1 U1004 ( .A1(n916), .A2(G401), .ZN(n913) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(n916), .ZN(G319) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1013 ( .A(G16), .B(KEYINPUT56), .Z(n943) );
  XNOR2_X1 U1014 ( .A(G1966), .B(G168), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(KEYINPUT57), .ZN(n929) );
  XNOR2_X1 U1017 ( .A(n920), .B(G1341), .ZN(n927) );
  XNOR2_X1 U1018 ( .A(G1961), .B(KEYINPUT118), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n921), .B(G301), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G1348), .B(n922), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT119), .B(n925), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n940) );
  NAND2_X1 U1025 ( .A1(G1971), .A2(G303), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n935) );
  XOR2_X1 U1027 ( .A(G1956), .B(G299), .Z(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(KEYINPUT120), .B(n938), .ZN(n939) );
  NOR2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1033 ( .A(KEYINPUT121), .B(n941), .Z(n942) );
  NOR2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n1025) );
  XOR2_X1 U1035 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n968) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(G1956), .B(G20), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n951) );
  XOR2_X1 U1039 ( .A(KEYINPUT122), .B(G4), .Z(n947) );
  XNOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(n947), .B(n946), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G1981), .B(G6), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(n952), .B(KEYINPUT60), .ZN(n962) );
  XOR2_X1 U1046 ( .A(G1971), .B(G22), .Z(n955) );
  XOR2_X1 U1047 ( .A(G24), .B(KEYINPUT124), .Z(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(G1986), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(G1976), .Z(n956) );
  XNOR2_X1 U1051 ( .A(G23), .B(n956), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT58), .B(n959), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT125), .B(n960), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G21), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G5), .B(G1961), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n968), .B(n967), .ZN(n970) );
  INV_X1 U1061 ( .A(G16), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n971), .ZN(n995) );
  XOR2_X1 U1064 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n992) );
  XNOR2_X1 U1065 ( .A(G2090), .B(G35), .ZN(n987) );
  XNOR2_X1 U1066 ( .A(G32), .B(n972), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(n973), .B(G27), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G26), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G33), .B(G2072), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(KEYINPUT116), .B(n980), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(G28), .ZN(n984) );
  XOR2_X1 U1075 ( .A(G25), .B(G1991), .Z(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT115), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT53), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1080 ( .A(G2084), .B(G34), .Z(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT54), .B(n988), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n992), .B(n991), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(G29), .A2(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1023) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT51), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1009) );
  XNOR2_X1 U1090 ( .A(G160), .B(G2084), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT113), .B(n1007), .Z(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1017) );
  XOR2_X1 U1096 ( .A(G2072), .B(n1010), .Z(n1012) );
  XOR2_X1 U1097 ( .A(G164), .B(G2078), .Z(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1013), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1018), .Z(n1019) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1019), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(KEYINPUT114), .B(n1020), .Z(n1021) );
  NAND2_X1 U1105 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1026), .Z(n1027) );
  XNOR2_X1 U1109 ( .A(KEYINPUT127), .B(n1027), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

