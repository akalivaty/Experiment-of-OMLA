

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752;

  XNOR2_X1 U379 ( .A(n462), .B(G469), .ZN(n596) );
  XNOR2_X1 U380 ( .A(G110), .B(n460), .ZN(n727) );
  INV_X1 U381 ( .A(KEYINPUT70), .ZN(n413) );
  XNOR2_X2 U382 ( .A(n359), .B(n416), .ZN(n721) );
  NAND2_X1 U383 ( .A1(n393), .A2(n396), .ZN(n359) );
  INV_X1 U384 ( .A(G953), .ZN(n737) );
  NOR2_X2 U385 ( .A1(G237), .A2(G953), .ZN(n450) );
  NOR2_X2 U386 ( .A1(n557), .A2(n690), .ZN(n559) );
  XNOR2_X2 U387 ( .A(n457), .B(G472), .ZN(n541) );
  XNOR2_X2 U388 ( .A(n464), .B(KEYINPUT20), .ZN(n477) );
  XNOR2_X2 U389 ( .A(n526), .B(n412), .ZN(n458) );
  XNOR2_X2 U390 ( .A(n413), .B(G131), .ZN(n526) );
  NOR2_X1 U391 ( .A1(n721), .A2(n736), .ZN(n665) );
  XOR2_X1 U392 ( .A(KEYINPUT6), .B(n687), .Z(n583) );
  INV_X2 U393 ( .A(n541), .ZN(n687) );
  NAND2_X1 U394 ( .A1(n665), .A2(KEYINPUT2), .ZN(n668) );
  NOR2_X1 U395 ( .A1(n585), .A2(n584), .ZN(n662) );
  XNOR2_X1 U396 ( .A(n392), .B(KEYINPUT19), .ZN(n597) );
  XNOR2_X1 U397 ( .A(n596), .B(KEYINPUT1), .ZN(n540) );
  OR2_X2 U398 ( .A1(n721), .A2(n388), .ZN(n628) );
  XNOR2_X2 U399 ( .A(n535), .B(n534), .ZN(n745) );
  XOR2_X2 U400 ( .A(n458), .B(n471), .Z(n733) );
  NOR2_X1 U401 ( .A1(n749), .A2(n748), .ZN(n406) );
  NOR2_X1 U402 ( .A1(n652), .A2(n752), .ZN(n551) );
  NOR2_X1 U403 ( .A1(G902), .A2(n708), .ZN(n462) );
  XNOR2_X1 U404 ( .A(n381), .B(n456), .ZN(n382) );
  XNOR2_X1 U405 ( .A(n458), .B(n410), .ZN(n456) );
  NAND2_X1 U406 ( .A1(n628), .A2(n627), .ZN(n640) );
  AND2_X2 U407 ( .A1(n640), .A2(n668), .ZN(n712) );
  XOR2_X1 U408 ( .A(KEYINPUT79), .B(KEYINPUT101), .Z(n452) );
  NOR2_X1 U409 ( .A1(n415), .A2(n750), .ZN(n414) );
  INV_X1 U410 ( .A(n664), .ZN(n415) );
  XNOR2_X1 U411 ( .A(n616), .B(KEYINPUT48), .ZN(n387) );
  AND2_X1 U412 ( .A1(n405), .A2(n377), .ZN(n616) );
  NOR2_X1 U413 ( .A1(n361), .A2(n615), .ZN(n377) );
  NOR2_X1 U414 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U415 ( .A1(n553), .A2(n552), .ZN(n399) );
  XNOR2_X1 U416 ( .A(n420), .B(G125), .ZN(n489) );
  INV_X1 U417 ( .A(G146), .ZN(n420) );
  NAND2_X1 U418 ( .A1(n446), .A2(n445), .ZN(n448) );
  XOR2_X1 U419 ( .A(G122), .B(G107), .Z(n508) );
  XNOR2_X1 U420 ( .A(G113), .B(G143), .ZN(n520) );
  BUF_X1 U421 ( .A(n540), .Z(n680) );
  XNOR2_X1 U422 ( .A(n373), .B(n502), .ZN(n503) );
  INV_X1 U423 ( .A(KEYINPUT0), .ZN(n502) );
  NAND2_X1 U424 ( .A1(n597), .A2(n501), .ZN(n373) );
  INV_X1 U425 ( .A(n670), .ZN(n409) );
  XNOR2_X1 U426 ( .A(n433), .B(n485), .ZN(n708) );
  XNOR2_X1 U427 ( .A(n436), .B(n459), .ZN(n435) );
  XNOR2_X1 U428 ( .A(n432), .B(n431), .ZN(n604) );
  INV_X1 U429 ( .A(KEYINPUT39), .ZN(n431) );
  AND2_X1 U430 ( .A1(n592), .A2(n364), .ZN(n422) );
  XNOR2_X1 U431 ( .A(n423), .B(n531), .ZN(n561) );
  OR2_X1 U432 ( .A1(n631), .A2(G902), .ZN(n423) );
  INV_X1 U433 ( .A(n557), .ZN(n554) );
  NAND2_X1 U434 ( .A1(n712), .A2(n368), .ZN(n428) );
  NOR2_X1 U435 ( .A1(n427), .A2(n716), .ZN(n426) );
  NAND2_X1 U436 ( .A1(n712), .A2(G469), .ZN(n386) );
  XNOR2_X1 U437 ( .A(n419), .B(n369), .ZN(n418) );
  XNOR2_X1 U438 ( .A(G116), .B(G113), .ZN(n440) );
  INV_X1 U439 ( .A(G128), .ZN(n444) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT104), .Z(n523) );
  XNOR2_X1 U441 ( .A(KEYINPUT12), .B(KEYINPUT103), .ZN(n522) );
  XOR2_X1 U442 ( .A(G104), .B(G122), .Z(n521) );
  XNOR2_X1 U443 ( .A(n400), .B(n489), .ZN(n491) );
  XNOR2_X1 U444 ( .A(n402), .B(n401), .ZN(n400) );
  XNOR2_X1 U445 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n402) );
  XNOR2_X1 U446 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n401) );
  NOR2_X1 U447 ( .A1(G902), .A2(G237), .ZN(n484) );
  XNOR2_X1 U448 ( .A(G146), .B(KEYINPUT78), .ZN(n451) );
  XNOR2_X1 U449 ( .A(KEYINPUT72), .B(G134), .ZN(n412) );
  XNOR2_X1 U450 ( .A(n449), .B(n411), .ZN(n410) );
  INV_X1 U451 ( .A(G137), .ZN(n411) );
  XNOR2_X1 U452 ( .A(n442), .B(n441), .ZN(n488) );
  XOR2_X1 U453 ( .A(KEYINPUT3), .B(G119), .Z(n441) );
  XNOR2_X1 U454 ( .A(n440), .B(n439), .ZN(n442) );
  INV_X1 U455 ( .A(KEYINPUT73), .ZN(n439) );
  NAND2_X1 U456 ( .A1(n387), .A2(n360), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n461), .B(KEYINPUT82), .ZN(n436) );
  XNOR2_X1 U458 ( .A(G146), .B(G140), .ZN(n461) );
  NAND2_X1 U459 ( .A1(n387), .A2(n414), .ZN(n736) );
  XNOR2_X1 U460 ( .A(n488), .B(n487), .ZN(n724) );
  XNOR2_X1 U461 ( .A(n486), .B(G122), .ZN(n487) );
  XOR2_X1 U462 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n486) );
  XOR2_X1 U463 ( .A(G107), .B(G104), .Z(n460) );
  INV_X1 U464 ( .A(KEYINPUT45), .ZN(n416) );
  XNOR2_X1 U465 ( .A(G119), .B(G128), .ZN(n467) );
  XNOR2_X1 U466 ( .A(G116), .B(G134), .ZN(n507) );
  XNOR2_X1 U467 ( .A(n528), .B(n424), .ZN(n631) );
  XNOR2_X1 U468 ( .A(n529), .B(n530), .ZN(n424) );
  XNOR2_X1 U469 ( .A(n403), .B(KEYINPUT22), .ZN(n547) );
  AND2_X1 U470 ( .A1(n539), .A2(n684), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n577), .B(KEYINPUT81), .ZN(n587) );
  NOR2_X1 U472 ( .A1(n575), .A2(n581), .ZN(n576) );
  XNOR2_X1 U473 ( .A(n372), .B(KEYINPUT28), .ZN(n595) );
  OR2_X1 U474 ( .A1(n593), .A2(n594), .ZN(n372) );
  NAND2_X1 U475 ( .A1(n379), .A2(n378), .ZN(n575) );
  INV_X1 U476 ( .A(n596), .ZN(n378) );
  INV_X1 U477 ( .A(n679), .ZN(n379) );
  XNOR2_X1 U478 ( .A(n603), .B(n421), .ZN(n645) );
  INV_X1 U479 ( .A(KEYINPUT114), .ZN(n421) );
  NOR2_X1 U480 ( .A1(n547), .A2(n618), .ZN(n567) );
  NOR2_X1 U481 ( .A1(n604), .A2(n603), .ZN(n606) );
  XNOR2_X1 U482 ( .A(n391), .B(n390), .ZN(n584) );
  INV_X1 U483 ( .A(KEYINPUT36), .ZN(n390) );
  NOR2_X1 U484 ( .A1(n617), .A2(n621), .ZN(n391) );
  NAND2_X1 U485 ( .A1(n428), .A2(n426), .ZN(n425) );
  INV_X1 U486 ( .A(KEYINPUT122), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n385), .A2(n430), .ZN(n384) );
  XNOR2_X1 U488 ( .A(n386), .B(n370), .ZN(n385) );
  NAND2_X1 U489 ( .A1(n418), .A2(n430), .ZN(n417) );
  AND2_X1 U490 ( .A1(n414), .A2(n623), .ZN(n360) );
  XOR2_X1 U491 ( .A(n614), .B(KEYINPUT76), .Z(n361) );
  INV_X1 U492 ( .A(n683), .ZN(n376) );
  XOR2_X1 U493 ( .A(KEYINPUT64), .B(KEYINPUT4), .Z(n362) );
  XOR2_X1 U494 ( .A(n489), .B(n469), .Z(n363) );
  AND2_X1 U495 ( .A1(n684), .A2(n670), .ZN(n364) );
  AND2_X1 U496 ( .A1(n645), .A2(n422), .ZN(n365) );
  XOR2_X1 U497 ( .A(n643), .B(n642), .Z(n366) );
  XOR2_X1 U498 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n367) );
  AND2_X1 U499 ( .A1(n366), .A2(G472), .ZN(n368) );
  XOR2_X1 U500 ( .A(n639), .B(n638), .Z(n369) );
  XOR2_X1 U501 ( .A(n708), .B(n707), .Z(n370) );
  XOR2_X1 U502 ( .A(n641), .B(KEYINPUT56), .Z(n371) );
  NOR2_X1 U503 ( .A1(n634), .A2(n716), .ZN(n374) );
  INV_X1 U504 ( .A(n716), .ZN(n430) );
  NAND2_X1 U505 ( .A1(n519), .A2(G210), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n450), .B(KEYINPUT80), .ZN(n519) );
  XNOR2_X1 U507 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U508 ( .A(n455), .B(n488), .ZN(n381) );
  XNOR2_X1 U509 ( .A(n374), .B(n636), .ZN(G60) );
  AND2_X1 U510 ( .A1(n567), .A2(n375), .ZN(n568) );
  NOR2_X1 U511 ( .A1(n583), .A2(n376), .ZN(n375) );
  NAND2_X1 U512 ( .A1(n629), .A2(n640), .ZN(n633) );
  XNOR2_X1 U513 ( .A(n727), .B(n435), .ZN(n434) );
  XNOR2_X1 U514 ( .A(n733), .B(n434), .ZN(n433) );
  XNOR2_X1 U515 ( .A(n480), .B(KEYINPUT97), .ZN(n481) );
  NAND2_X1 U516 ( .A1(n395), .A2(KEYINPUT66), .ZN(n394) );
  XNOR2_X1 U517 ( .A(n380), .B(n367), .ZN(n669) );
  NAND2_X1 U518 ( .A1(n583), .A2(n483), .ZN(n380) );
  XNOR2_X1 U519 ( .A(n485), .B(n382), .ZN(n643) );
  XNOR2_X2 U520 ( .A(n734), .B(G101), .ZN(n485) );
  XNOR2_X2 U521 ( .A(n506), .B(n362), .ZN(n734) );
  XNOR2_X1 U522 ( .A(n384), .B(n383), .ZN(G54) );
  NAND2_X1 U523 ( .A1(n583), .A2(n365), .ZN(n617) );
  NAND2_X1 U524 ( .A1(n580), .A2(n670), .ZN(n392) );
  XNOR2_X2 U525 ( .A(n496), .B(n437), .ZN(n580) );
  NAND2_X1 U526 ( .A1(n394), .A2(n551), .ZN(n393) );
  NAND2_X1 U527 ( .A1(n538), .A2(n537), .ZN(n395) );
  AND2_X1 U528 ( .A1(n397), .A2(n399), .ZN(n396) );
  NOR2_X1 U529 ( .A1(n570), .A2(n398), .ZN(n397) );
  NAND2_X1 U530 ( .A1(n744), .A2(n569), .ZN(n398) );
  INV_X1 U531 ( .A(n503), .ZN(n557) );
  NAND2_X1 U532 ( .A1(n503), .A2(n404), .ZN(n403) );
  XNOR2_X1 U533 ( .A(n406), .B(n611), .ZN(n405) );
  NAND2_X1 U534 ( .A1(n576), .A2(n407), .ZN(n577) );
  XNOR2_X1 U535 ( .A(n408), .B(KEYINPUT30), .ZN(n407) );
  NOR2_X1 U536 ( .A1(n541), .A2(n409), .ZN(n408) );
  XNOR2_X1 U537 ( .A(n724), .B(n492), .ZN(n493) );
  XNOR2_X1 U538 ( .A(n494), .B(n493), .ZN(n637) );
  XNOR2_X1 U539 ( .A(n417), .B(n371), .ZN(G51) );
  NAND2_X1 U540 ( .A1(n712), .A2(G210), .ZN(n419) );
  NOR2_X1 U541 ( .A1(n429), .A2(n425), .ZN(n644) );
  NOR2_X1 U542 ( .A1(n366), .A2(G472), .ZN(n427) );
  NOR2_X1 U543 ( .A1(n712), .A2(n366), .ZN(n429) );
  NAND2_X1 U544 ( .A1(n587), .A2(n671), .ZN(n432) );
  NOR2_X2 U545 ( .A1(n533), .A2(n586), .ZN(n535) );
  AND2_X1 U546 ( .A1(n495), .A2(G210), .ZN(n437) );
  INV_X1 U547 ( .A(KEYINPUT68), .ZN(n536) );
  INV_X1 U548 ( .A(G143), .ZN(n447) );
  XNOR2_X1 U549 ( .A(n454), .B(n453), .ZN(n455) );
  INV_X1 U550 ( .A(KEYINPUT59), .ZN(n630) );
  XNOR2_X1 U551 ( .A(n631), .B(n630), .ZN(n632) );
  INV_X1 U552 ( .A(KEYINPUT123), .ZN(n635) );
  XNOR2_X1 U553 ( .A(n635), .B(KEYINPUT60), .ZN(n636) );
  NOR2_X1 U554 ( .A1(G952), .A2(n737), .ZN(n438) );
  XNOR2_X1 U555 ( .A(KEYINPUT94), .B(n438), .ZN(n716) );
  INV_X1 U556 ( .A(KEYINPUT65), .ZN(n443) );
  NAND2_X1 U557 ( .A1(G128), .A2(n443), .ZN(n446) );
  NAND2_X1 U558 ( .A1(n444), .A2(KEYINPUT65), .ZN(n445) );
  XNOR2_X2 U559 ( .A(n448), .B(n447), .ZN(n506) );
  XNOR2_X1 U560 ( .A(KEYINPUT5), .B(KEYINPUT100), .ZN(n449) );
  XNOR2_X1 U561 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U562 ( .A1(G902), .A2(n643), .ZN(n457) );
  XOR2_X1 U563 ( .A(G137), .B(KEYINPUT71), .Z(n471) );
  NAND2_X1 U564 ( .A1(G227), .A2(n737), .ZN(n459) );
  XOR2_X1 U565 ( .A(KEYINPUT21), .B(KEYINPUT99), .Z(n466) );
  XNOR2_X2 U566 ( .A(G902), .B(KEYINPUT15), .ZN(n463) );
  XOR2_X2 U567 ( .A(n463), .B(KEYINPUT95), .Z(n624) );
  NAND2_X1 U568 ( .A1(G234), .A2(n624), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n477), .A2(G221), .ZN(n465) );
  XOR2_X1 U570 ( .A(n466), .B(n465), .Z(n684) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(G110), .Z(n468) );
  XNOR2_X1 U572 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U573 ( .A(KEYINPUT10), .B(G140), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n470), .B(n363), .ZN(n476) );
  XOR2_X1 U575 ( .A(n471), .B(KEYINPUT24), .Z(n474) );
  NAND2_X1 U576 ( .A1(G234), .A2(n737), .ZN(n472) );
  XOR2_X1 U577 ( .A(KEYINPUT8), .B(n472), .Z(n511) );
  NAND2_X1 U578 ( .A1(G221), .A2(n511), .ZN(n473) );
  XNOR2_X1 U579 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n476), .B(n475), .ZN(n714) );
  NOR2_X1 U581 ( .A1(n714), .A2(G902), .ZN(n482) );
  XOR2_X1 U582 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n479) );
  NAND2_X1 U583 ( .A1(n477), .A2(G217), .ZN(n478) );
  XNOR2_X1 U584 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X2 U585 ( .A(n482), .B(n481), .ZN(n582) );
  NAND2_X1 U586 ( .A1(n684), .A2(n582), .ZN(n679) );
  NOR2_X2 U587 ( .A1(n540), .A2(n679), .ZN(n556) );
  XNOR2_X1 U588 ( .A(n556), .B(KEYINPUT112), .ZN(n483) );
  INV_X1 U589 ( .A(n669), .ZN(n504) );
  XNOR2_X1 U590 ( .A(n484), .B(KEYINPUT77), .ZN(n495) );
  NAND2_X1 U591 ( .A1(G214), .A2(n495), .ZN(n670) );
  XNOR2_X1 U592 ( .A(n727), .B(n485), .ZN(n494) );
  NAND2_X1 U593 ( .A1(G224), .A2(n737), .ZN(n490) );
  XOR2_X1 U594 ( .A(n491), .B(n490), .Z(n492) );
  NAND2_X1 U595 ( .A1(n637), .A2(n624), .ZN(n496) );
  NAND2_X1 U596 ( .A1(G234), .A2(G237), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n497), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U598 ( .A1(G952), .A2(n498), .ZN(n698) );
  NOR2_X1 U599 ( .A1(G953), .A2(n698), .ZN(n574) );
  NAND2_X1 U600 ( .A1(G902), .A2(n498), .ZN(n571) );
  INV_X1 U601 ( .A(G898), .ZN(n719) );
  NAND2_X1 U602 ( .A1(G953), .A2(n719), .ZN(n728) );
  NOR2_X1 U603 ( .A1(n571), .A2(n728), .ZN(n499) );
  NOR2_X1 U604 ( .A1(n574), .A2(n499), .ZN(n500) );
  XOR2_X1 U605 ( .A(KEYINPUT96), .B(n500), .Z(n501) );
  NAND2_X1 U606 ( .A1(n504), .A2(n554), .ZN(n505) );
  XNOR2_X1 U607 ( .A(n505), .B(KEYINPUT34), .ZN(n533) );
  INV_X1 U608 ( .A(n506), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n510), .B(n509), .ZN(n513) );
  NAND2_X1 U611 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U612 ( .A(n513), .B(n512), .ZN(n515) );
  XOR2_X1 U613 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n514) );
  XNOR2_X1 U614 ( .A(n515), .B(n514), .ZN(n710) );
  NOR2_X1 U615 ( .A1(G902), .A2(n710), .ZN(n516) );
  XNOR2_X1 U616 ( .A(G478), .B(n516), .ZN(n560) );
  XOR2_X1 U617 ( .A(KEYINPUT13), .B(KEYINPUT106), .Z(n518) );
  XNOR2_X1 U618 ( .A(KEYINPUT107), .B(G475), .ZN(n517) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n531) );
  NAND2_X1 U620 ( .A1(n519), .A2(G214), .ZN(n530) );
  XNOR2_X1 U621 ( .A(n521), .B(n520), .ZN(n525) );
  XNOR2_X1 U622 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U623 ( .A(n525), .B(n524), .ZN(n529) );
  XNOR2_X1 U624 ( .A(n526), .B(KEYINPUT105), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n527), .B(n363), .ZN(n528) );
  NOR2_X1 U626 ( .A1(n560), .A2(n561), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT113), .ZN(n586) );
  INV_X1 U628 ( .A(KEYINPUT35), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n745), .B(n536), .ZN(n538) );
  INV_X1 U630 ( .A(KEYINPUT44), .ZN(n537) );
  INV_X1 U631 ( .A(n684), .ZN(n594) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n673) );
  INV_X1 U633 ( .A(n673), .ZN(n539) );
  INV_X1 U634 ( .A(n680), .ZN(n618) );
  NAND2_X1 U635 ( .A1(n567), .A2(n541), .ZN(n542) );
  NOR2_X1 U636 ( .A1(n582), .A2(n542), .ZN(n652) );
  INV_X1 U637 ( .A(KEYINPUT32), .ZN(n550) );
  INV_X1 U638 ( .A(n583), .ZN(n543) );
  XOR2_X1 U639 ( .A(KEYINPUT85), .B(n543), .Z(n545) );
  XOR2_X1 U640 ( .A(KEYINPUT93), .B(n680), .Z(n585) );
  INV_X1 U641 ( .A(n585), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U643 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U644 ( .A(n582), .B(KEYINPUT110), .ZN(n683) );
  NAND2_X1 U645 ( .A1(n548), .A2(n376), .ZN(n549) );
  XNOR2_X1 U646 ( .A(n550), .B(n549), .ZN(n752) );
  NAND2_X1 U647 ( .A1(KEYINPUT68), .A2(n551), .ZN(n553) );
  AND2_X1 U648 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n552) );
  NOR2_X1 U649 ( .A1(n687), .A2(n575), .ZN(n555) );
  NAND2_X1 U650 ( .A1(n555), .A2(n554), .ZN(n648) );
  NAND2_X1 U651 ( .A1(n687), .A2(n556), .ZN(n690) );
  XNOR2_X1 U652 ( .A(KEYINPUT31), .B(KEYINPUT102), .ZN(n558) );
  XNOR2_X1 U653 ( .A(n559), .B(n558), .ZN(n660) );
  NAND2_X1 U654 ( .A1(n648), .A2(n660), .ZN(n563) );
  INV_X1 U655 ( .A(n560), .ZN(n562) );
  OR2_X1 U656 ( .A1(n562), .A2(n561), .ZN(n603) );
  NAND2_X1 U657 ( .A1(n562), .A2(n561), .ZN(n659) );
  XNOR2_X1 U658 ( .A(KEYINPUT108), .B(n659), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n603), .A2(n578), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n563), .A2(n590), .ZN(n564) );
  XNOR2_X1 U661 ( .A(n564), .B(KEYINPUT109), .ZN(n566) );
  NOR2_X1 U662 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n568), .B(KEYINPUT111), .ZN(n744) );
  AND2_X1 U664 ( .A1(KEYINPUT44), .A2(n745), .ZN(n570) );
  OR2_X1 U665 ( .A1(n737), .A2(n571), .ZN(n572) );
  NOR2_X1 U666 ( .A1(G900), .A2(n572), .ZN(n573) );
  NOR2_X1 U667 ( .A1(n574), .A2(n573), .ZN(n581) );
  XOR2_X1 U668 ( .A(KEYINPUT38), .B(n580), .Z(n671) );
  NOR2_X1 U669 ( .A1(n578), .A2(n604), .ZN(n579) );
  XNOR2_X1 U670 ( .A(KEYINPUT118), .B(n579), .ZN(n750) );
  INV_X1 U671 ( .A(n580), .ZN(n621) );
  NOR2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n592) );
  XNOR2_X1 U673 ( .A(KEYINPUT91), .B(n662), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n621), .A2(n586), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U676 ( .A(KEYINPUT116), .B(n589), .Z(n751) );
  INV_X1 U677 ( .A(n590), .ZN(n675) );
  NAND2_X1 U678 ( .A1(n675), .A2(KEYINPUT47), .ZN(n591) );
  XOR2_X1 U679 ( .A(n591), .B(KEYINPUT87), .Z(n599) );
  NAND2_X1 U680 ( .A1(n687), .A2(n592), .ZN(n593) );
  NOR2_X1 U681 ( .A1(n596), .A2(n595), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n607), .A2(n597), .ZN(n655) );
  NAND2_X1 U683 ( .A1(n655), .A2(KEYINPUT47), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U685 ( .A1(n751), .A2(n600), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n615) );
  XOR2_X1 U687 ( .A(KEYINPUT117), .B(KEYINPUT40), .Z(n605) );
  XNOR2_X1 U688 ( .A(n606), .B(n605), .ZN(n749) );
  INV_X1 U689 ( .A(n607), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n671), .A2(n670), .ZN(n674) );
  NOR2_X1 U691 ( .A1(n674), .A2(n673), .ZN(n608) );
  XNOR2_X1 U692 ( .A(n608), .B(KEYINPUT41), .ZN(n699) );
  NOR2_X1 U693 ( .A1(n609), .A2(n699), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n610), .B(KEYINPUT42), .ZN(n748) );
  XNOR2_X1 U695 ( .A(KEYINPUT46), .B(KEYINPUT90), .ZN(n611) );
  XNOR2_X1 U696 ( .A(KEYINPUT69), .B(KEYINPUT47), .ZN(n613) );
  NOR2_X1 U697 ( .A1(n675), .A2(n655), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U700 ( .A(KEYINPUT115), .B(KEYINPUT43), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n664) );
  AND2_X1 U703 ( .A1(n668), .A2(G475), .ZN(n629) );
  INV_X1 U704 ( .A(n624), .ZN(n623) );
  XOR2_X1 U705 ( .A(n624), .B(KEYINPUT88), .Z(n625) );
  NAND2_X1 U706 ( .A1(n625), .A2(KEYINPUT2), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT67), .B(n626), .Z(n627) );
  XNOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n637), .B(KEYINPUT92), .ZN(n638) );
  INV_X1 U710 ( .A(KEYINPUT89), .ZN(n641) );
  XOR2_X1 U711 ( .A(KEYINPUT119), .B(KEYINPUT62), .Z(n642) );
  XOR2_X1 U712 ( .A(KEYINPUT63), .B(n644), .Z(G57) );
  INV_X1 U713 ( .A(n645), .ZN(n657) );
  NOR2_X1 U714 ( .A1(n657), .A2(n648), .ZN(n646) );
  XOR2_X1 U715 ( .A(KEYINPUT120), .B(n646), .Z(n647) );
  XNOR2_X1 U716 ( .A(G104), .B(n647), .ZN(G6) );
  NOR2_X1 U717 ( .A1(n659), .A2(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U720 ( .A(G107), .B(n651), .ZN(G9) );
  XOR2_X1 U721 ( .A(G110), .B(n652), .Z(G12) );
  NOR2_X1 U722 ( .A1(n659), .A2(n655), .ZN(n654) );
  XNOR2_X1 U723 ( .A(G128), .B(KEYINPUT29), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(G30) );
  NOR2_X1 U725 ( .A1(n657), .A2(n655), .ZN(n656) );
  XOR2_X1 U726 ( .A(G146), .B(n656), .Z(G48) );
  NOR2_X1 U727 ( .A1(n657), .A2(n660), .ZN(n658) );
  XOR2_X1 U728 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U730 ( .A(G116), .B(n661), .Z(G18) );
  XNOR2_X1 U731 ( .A(G125), .B(n662), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U733 ( .A(G140), .B(n664), .ZN(G42) );
  NOR2_X1 U734 ( .A1(n665), .A2(KEYINPUT2), .ZN(n666) );
  XOR2_X1 U735 ( .A(KEYINPUT86), .B(n666), .Z(n667) );
  NAND2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n704) );
  BUF_X1 U737 ( .A(n669), .Z(n700) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n700), .A2(n678), .ZN(n695) );
  AND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U744 ( .A(n681), .B(KEYINPUT50), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n682), .B(KEYINPUT121), .ZN(n689) );
  NOR2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U747 ( .A(KEYINPUT49), .B(n685), .Z(n686) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U749 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U751 ( .A(KEYINPUT51), .B(n692), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n699), .A2(n693), .ZN(n694) );
  NOR2_X1 U753 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U754 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U761 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n707) );
  NAND2_X1 U762 ( .A1(G478), .A2(n712), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n716), .A2(n711), .ZN(G63) );
  NAND2_X1 U765 ( .A1(G217), .A2(n712), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(G66) );
  XOR2_X1 U768 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n718) );
  NAND2_X1 U769 ( .A1(G224), .A2(G953), .ZN(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U772 ( .A1(G953), .A2(n721), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n732) );
  XNOR2_X1 U774 ( .A(n724), .B(G101), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n725), .B(KEYINPUT125), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U778 ( .A(n730), .B(KEYINPUT126), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n732), .B(n731), .ZN(G69) );
  XOR2_X1 U780 ( .A(n734), .B(n733), .Z(n735) );
  XNOR2_X1 U781 ( .A(n363), .B(n735), .ZN(n739) );
  XNOR2_X1 U782 ( .A(n739), .B(n736), .ZN(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(n737), .ZN(n743) );
  XNOR2_X1 U784 ( .A(G227), .B(n739), .ZN(n740) );
  NAND2_X1 U785 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U786 ( .A1(G953), .A2(n741), .ZN(n742) );
  NAND2_X1 U787 ( .A1(n743), .A2(n742), .ZN(G72) );
  XNOR2_X1 U788 ( .A(n744), .B(G101), .ZN(G3) );
  INV_X1 U789 ( .A(n745), .ZN(n746) );
  XOR2_X1 U790 ( .A(G122), .B(n746), .Z(n747) );
  XNOR2_X1 U791 ( .A(n747), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U792 ( .A(G137), .B(n748), .Z(G39) );
  XOR2_X1 U793 ( .A(G131), .B(n749), .Z(G33) );
  XOR2_X1 U794 ( .A(G134), .B(n750), .Z(G36) );
  XOR2_X1 U795 ( .A(G143), .B(n751), .Z(G45) );
  XOR2_X1 U796 ( .A(G119), .B(n752), .Z(G21) );
endmodule

