

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  NOR2_X1 U327 ( .A1(n534), .A2(n459), .ZN(n574) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  INV_X1 U329 ( .A(KEYINPUT46), .ZN(n405) );
  XNOR2_X1 U330 ( .A(n438), .B(n295), .ZN(n371) );
  XNOR2_X1 U331 ( .A(n391), .B(n371), .ZN(n372) );
  INV_X1 U332 ( .A(KEYINPUT76), .ZN(n378) );
  XNOR2_X1 U333 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U334 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U335 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U336 ( .A(n381), .B(n380), .ZN(n383) );
  INV_X1 U337 ( .A(G211GAT), .ZN(n452) );
  INV_X1 U338 ( .A(G190GAT), .ZN(n460) );
  XOR2_X1 U339 ( .A(n347), .B(n346), .Z(n534) );
  XNOR2_X1 U340 ( .A(n452), .B(KEYINPUT126), .ZN(n453) );
  XNOR2_X1 U341 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(G1354GAT) );
  XNOR2_X1 U343 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(G8GAT), .B(G183GAT), .Z(n413) );
  XNOR2_X1 U345 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n399) );
  XNOR2_X1 U346 ( .A(n413), .B(n399), .ZN(n297) );
  XOR2_X1 U347 ( .A(G15GAT), .B(KEYINPUT70), .Z(n360) );
  XOR2_X1 U348 ( .A(G22GAT), .B(G155GAT), .Z(n325) );
  XNOR2_X1 U349 ( .A(n360), .B(n325), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n310) );
  XOR2_X1 U351 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n299) );
  NAND2_X1 U352 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(n300), .B(KEYINPUT12), .Z(n308) );
  XOR2_X1 U355 ( .A(G211GAT), .B(G78GAT), .Z(n302) );
  XNOR2_X1 U356 ( .A(G127GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U358 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n304) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(G64GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U363 ( .A(n310), .B(n309), .Z(n573) );
  INV_X1 U364 ( .A(n573), .ZN(n494) );
  XOR2_X1 U365 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n312) );
  XNOR2_X1 U366 ( .A(G218GAT), .B(G106GAT), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n329) );
  XOR2_X1 U368 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n314) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(n315), .B(KEYINPUT24), .Z(n321) );
  XOR2_X1 U372 ( .A(G78GAT), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U373 ( .A(KEYINPUT72), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n390) );
  XOR2_X1 U375 ( .A(KEYINPUT3), .B(KEYINPUT88), .Z(n319) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n447) );
  XNOR2_X1 U378 ( .A(n390), .B(n447), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n324) );
  XOR2_X1 U380 ( .A(G211GAT), .B(KEYINPUT21), .Z(n323) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n419) );
  XOR2_X1 U383 ( .A(n324), .B(n419), .Z(n327) );
  XOR2_X1 U384 ( .A(G50GAT), .B(G162GAT), .Z(n377) );
  XNOR2_X1 U385 ( .A(n377), .B(n325), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U387 ( .A(n329), .B(n328), .Z(n474) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G71GAT), .Z(n396) );
  XOR2_X1 U389 ( .A(G134GAT), .B(G99GAT), .Z(n331) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n396), .B(n332), .Z(n334) );
  NAND2_X1 U393 ( .A1(G227GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U395 ( .A(G176GAT), .B(KEYINPUT83), .Z(n336) );
  XNOR2_X1 U396 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U398 ( .A(G183GAT), .B(KEYINPUT84), .Z(n338) );
  XNOR2_X1 U399 ( .A(G15GAT), .B(KEYINPUT85), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U401 ( .A(n340), .B(n339), .Z(n345) );
  XNOR2_X1 U402 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n341) );
  XOR2_X1 U403 ( .A(n341), .B(KEYINPUT82), .Z(n448) );
  XOR2_X1 U404 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n343) );
  XNOR2_X1 U405 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n425) );
  XOR2_X1 U407 ( .A(n448), .B(n425), .Z(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U409 ( .A1(n474), .A2(n534), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n348), .B(KEYINPUT26), .ZN(n554) );
  XOR2_X1 U411 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n350) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(G29GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U414 ( .A(KEYINPUT69), .B(n351), .ZN(n382) );
  XOR2_X1 U415 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n353) );
  XNOR2_X1 U416 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n367) );
  XOR2_X1 U418 ( .A(G141GAT), .B(G22GAT), .Z(n355) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G50GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U421 ( .A(KEYINPUT67), .B(G8GAT), .Z(n357) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(G197GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U425 ( .A(G113GAT), .B(G1GAT), .Z(n439) );
  XOR2_X1 U426 ( .A(n360), .B(KEYINPUT29), .Z(n362) );
  NAND2_X1 U427 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n439), .B(n363), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U431 ( .A(n367), .B(n366), .Z(n368) );
  XNOR2_X1 U432 ( .A(n382), .B(n368), .ZN(n577) );
  INV_X1 U433 ( .A(n577), .ZN(n567) );
  INV_X1 U434 ( .A(KEYINPUT78), .ZN(n384) );
  XOR2_X1 U435 ( .A(G92GAT), .B(G85GAT), .Z(n370) );
  XNOR2_X1 U436 ( .A(G99GAT), .B(G106GAT), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n391) );
  XOR2_X1 U438 ( .A(G134GAT), .B(KEYINPUT75), .Z(n438) );
  XOR2_X1 U439 ( .A(n372), .B(KEYINPUT10), .Z(n376) );
  XOR2_X1 U440 ( .A(KEYINPUT77), .B(G218GAT), .Z(n374) );
  XNOR2_X1 U441 ( .A(G36GAT), .B(G190GAT), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n417) );
  XNOR2_X1 U443 ( .A(n417), .B(KEYINPUT9), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n377), .B(KEYINPUT11), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n403) );
  XNOR2_X1 U447 ( .A(n384), .B(n403), .ZN(n548) );
  XOR2_X1 U448 ( .A(KEYINPUT36), .B(n548), .Z(n587) );
  NOR2_X1 U449 ( .A1(n494), .A2(n587), .ZN(n386) );
  XOR2_X1 U450 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n401) );
  XOR2_X1 U452 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n388) );
  NAND2_X1 U453 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U455 ( .A(n389), .B(KEYINPUT32), .Z(n393) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(G176GAT), .B(G64GAT), .Z(n414) );
  XOR2_X1 U459 ( .A(n394), .B(n414), .Z(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n395) );
  XOR2_X1 U461 ( .A(n400), .B(n399), .Z(n582) );
  NAND2_X1 U462 ( .A1(n401), .A2(n582), .ZN(n402) );
  NOR2_X1 U463 ( .A1(n567), .A2(n402), .ZN(n411) );
  XNOR2_X1 U464 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n404) );
  XOR2_X1 U465 ( .A(n404), .B(n582), .Z(n556) );
  OR2_X1 U466 ( .A1(n556), .A2(n577), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n407) );
  NOR2_X1 U468 ( .A1(n573), .A2(n407), .ZN(n408) );
  NAND2_X1 U469 ( .A1(n403), .A2(n408), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n409), .B(KEYINPUT47), .ZN(n410) );
  NOR2_X1 U471 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n412), .B(KEYINPUT48), .ZN(n531) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n423) );
  XOR2_X1 U474 ( .A(G92GAT), .B(KEYINPUT94), .Z(n416) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U477 ( .A(n418), .B(n417), .Z(n421) );
  XNOR2_X1 U478 ( .A(G204GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n523) );
  NOR2_X1 U482 ( .A1(n531), .A2(n523), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n426), .B(KEYINPUT54), .ZN(n457) );
  XOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n428) );
  XNOR2_X1 U485 ( .A(G120GAT), .B(G155GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U487 ( .A(KEYINPUT5), .B(G57GAT), .Z(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n432), .B(n431), .Z(n437) );
  XOR2_X1 U491 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n434) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(KEYINPUT93), .B(n435), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U496 ( .A(n438), .B(G162GAT), .Z(n441) );
  XNOR2_X1 U497 ( .A(n439), .B(G148GAT), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U500 ( .A(G29GAT), .B(G85GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n521) );
  NAND2_X1 U504 ( .A1(n457), .A2(n521), .ZN(n450) );
  NOR2_X1 U505 ( .A1(n554), .A2(n450), .ZN(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT123), .B(n451), .ZN(n586) );
  NOR2_X1 U507 ( .A1(n494), .A2(n586), .ZN(n454) );
  INV_X1 U508 ( .A(n474), .ZN(n455) );
  AND2_X1 U509 ( .A1(n521), .A2(n455), .ZN(n456) );
  AND2_X1 U510 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT55), .ZN(n459) );
  NAND2_X1 U512 ( .A1(n574), .A2(n548), .ZN(n463) );
  XOR2_X1 U513 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n461) );
  XOR2_X1 U514 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n465) );
  XNOR2_X1 U515 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n465), .B(n464), .ZN(n483) );
  AND2_X1 U517 ( .A1(n567), .A2(n582), .ZN(n498) );
  NOR2_X1 U518 ( .A1(n534), .A2(n523), .ZN(n466) );
  NOR2_X1 U519 ( .A1(n474), .A2(n466), .ZN(n467) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n467), .Z(n470) );
  XOR2_X1 U521 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n468) );
  XNOR2_X1 U522 ( .A(n523), .B(n468), .ZN(n475) );
  NOR2_X1 U523 ( .A1(n554), .A2(n475), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U525 ( .A(KEYINPUT96), .B(n471), .Z(n472) );
  NAND2_X1 U526 ( .A1(n472), .A2(n521), .ZN(n473) );
  XNOR2_X1 U527 ( .A(n473), .B(KEYINPUT97), .ZN(n478) );
  XNOR2_X1 U528 ( .A(n474), .B(KEYINPUT28), .ZN(n537) );
  NOR2_X1 U529 ( .A1(n475), .A2(n521), .ZN(n532) );
  NAND2_X1 U530 ( .A1(n534), .A2(n532), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n537), .A2(n476), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n478), .A2(n477), .ZN(n492) );
  XOR2_X1 U533 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n480) );
  OR2_X1 U534 ( .A1(n494), .A2(n548), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n480), .B(n479), .ZN(n481) );
  NOR2_X1 U536 ( .A1(n492), .A2(n481), .ZN(n509) );
  NAND2_X1 U537 ( .A1(n498), .A2(n509), .ZN(n489) );
  NOR2_X1 U538 ( .A1(n521), .A2(n489), .ZN(n482) );
  XOR2_X1 U539 ( .A(n483), .B(n482), .Z(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT98), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n523), .A2(n489), .ZN(n485) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n534), .A2(n489), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  INV_X1 U547 ( .A(n537), .ZN(n527) );
  NOR2_X1 U548 ( .A1(n527), .A2(n489), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(n490), .Z(n491) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(KEYINPUT105), .Z(n500) );
  NOR2_X1 U552 ( .A1(n587), .A2(n492), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n494), .A2(n493), .ZN(n497) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT37), .Z(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT103), .B(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n519) );
  NAND2_X1 U557 ( .A1(n498), .A2(n519), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n500), .B(n499), .ZN(n507) );
  NOR2_X1 U559 ( .A1(n507), .A2(n521), .ZN(n502) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n507), .A2(n523), .ZN(n503) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  XNOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n505) );
  NOR2_X1 U565 ( .A1(n534), .A2(n507), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U567 ( .A(G43GAT), .B(n506), .Z(G1330GAT) );
  NOR2_X1 U568 ( .A1(n527), .A2(n507), .ZN(n508) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(n556), .Z(n569) );
  AND2_X1 U571 ( .A1(n569), .A2(n577), .ZN(n520) );
  NAND2_X1 U572 ( .A1(n520), .A2(n509), .ZN(n516) );
  NOR2_X1 U573 ( .A1(n521), .A2(n516), .ZN(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n516), .ZN(n513) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n534), .A2(n516), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n527), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n521), .A2(n526), .ZN(n522) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n534), .A2(n526), .ZN(n525) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  INV_X1 U596 ( .A(n531), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n553) );
  NOR2_X1 U598 ( .A1(n534), .A2(n553), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT111), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n567), .A2(n549), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n540) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT112), .B(n541), .Z(n543) );
  NAND2_X1 U607 ( .A1(n549), .A2(n569), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n545) );
  NAND2_X1 U611 ( .A1(n549), .A2(n573), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NOR2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n562), .A2(n567), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  INV_X1 U621 ( .A(n562), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n556), .A2(n565), .ZN(n558) );
  XNOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(n559), .B(KEYINPUT52), .Z(n561) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n573), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NOR2_X1 U631 ( .A1(n403), .A2(n565), .ZN(n566) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n574), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n571) );
  NAND2_X1 U636 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(n572), .ZN(G1349GAT) );
  XOR2_X1 U639 ( .A(G183GAT), .B(KEYINPUT121), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n586), .ZN(n581) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT60), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n586), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n585), .B(G204GAT), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

