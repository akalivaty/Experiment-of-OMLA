//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT68), .B1(new_n188), .B2(G119), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(G116), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n191), .B(new_n192), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n202), .A2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n200), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n198), .A2(new_n206), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n199), .A2(new_n201), .A3(new_n203), .A4(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(G137), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n216), .B2(G137), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(KEYINPUT64), .A3(KEYINPUT11), .A4(G134), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(G134), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n218), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n213), .A2(new_n223), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n214), .A2(new_n215), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n220), .A2(new_n222), .A3(new_n231), .A4(new_n224), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT65), .A2(G131), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n217), .A2(new_n233), .A3(new_n220), .A4(new_n222), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT0), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(new_n198), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT0), .B(G128), .Z(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT30), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n230), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n230), .B2(new_n243), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n197), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n196), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n195), .B(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n230), .A3(new_n243), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n253), .B(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n250), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n249), .B1(new_n243), .B2(new_n230), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT28), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n187), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  OAI21_X1  g081(.A(G472), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(G472), .A2(G902), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n250), .A2(new_n256), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n250), .A2(new_n273), .A3(new_n256), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n247), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT71), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n247), .A3(new_n274), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT31), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n260), .A2(new_n262), .ZN(new_n280));
  INV_X1    g094(.A(new_n256), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT32), .B(new_n269), .C1(new_n279), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n276), .A2(new_n278), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n288), .B(new_n282), .C1(new_n283), .C2(new_n278), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT32), .B1(new_n289), .B2(new_n269), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n269), .B1(new_n279), .B2(new_n284), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n268), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT84), .Z(new_n297));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n298));
  INV_X1    g112(.A(G107), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(G104), .ZN(new_n300));
  INV_X1    g114(.A(G104), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT80), .A3(G107), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n301), .A2(G107), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT3), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND4_X1   g120(.A1(new_n305), .A2(new_n299), .A3(KEYINPUT3), .A4(G104), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G101), .ZN(new_n309));
  INV_X1    g123(.A(G101), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n310), .B(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(KEYINPUT4), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n313), .A3(G101), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n197), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n299), .A2(G104), .ZN(new_n316));
  OAI21_X1  g130(.A(G101), .B1(new_n304), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n195), .A2(new_n196), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n189), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(G113), .B(new_n322), .C1(new_n195), .C2(new_n321), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G110), .B(G122), .Z(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n315), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(KEYINPUT6), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n242), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n205), .A2(new_n210), .A3(new_n212), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G953), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G224), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n335), .B(new_n337), .Z(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n325), .A2(new_n339), .A3(new_n326), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n330), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT7), .A4(new_n337), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT88), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT87), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(KEYINPUT7), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n344), .B(new_n345), .C1(KEYINPUT87), .C2(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n323), .A2(new_n320), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n317), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n326), .B(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n343), .A2(new_n346), .A3(new_n329), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n354), .A3(new_n187), .ZN(new_n355));
  OAI21_X1  g169(.A(G210), .B1(G237), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n341), .A2(new_n354), .A3(new_n187), .A4(new_n356), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n297), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT93), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n331), .A2(KEYINPUT16), .A3(G140), .ZN(new_n362));
  XNOR2_X1  g176(.A(G125), .B(G140), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(KEYINPUT16), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G146), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(G146), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n254), .A2(G143), .A3(G214), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(G143), .B1(new_n254), .B2(G214), .ZN(new_n371));
  OAI21_X1  g185(.A(G131), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT17), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(KEYINPUT16), .ZN(new_n375));
  INV_X1    g189(.A(new_n362), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n200), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT93), .A3(new_n365), .ZN(new_n379));
  INV_X1    g193(.A(G237), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n336), .A3(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n202), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n218), .A3(new_n369), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n372), .A2(new_n373), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n368), .A2(new_n374), .A3(new_n379), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(KEYINPUT89), .A3(new_n369), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT18), .A2(G131), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n363), .B(new_n200), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(G113), .B(G122), .Z(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT92), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(new_n301), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(G104), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n372), .A2(new_n383), .B1(G146), .B2(new_n364), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n363), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT19), .B1(new_n363), .B2(KEYINPUT90), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n200), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n388), .A2(new_n389), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n401), .B2(KEYINPUT91), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n400), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n390), .A2(KEYINPUT91), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n394), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G475), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n187), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT20), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n405), .A2(new_n409), .A3(new_n406), .A4(new_n187), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n385), .A2(new_n390), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n395), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n394), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n406), .B1(new_n414), .B2(new_n187), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT96), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n187), .B(new_n336), .C1(G234), .C2(G237), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G952), .ZN(new_n423));
  AOI211_X1 g237(.A(G953), .B(new_n423), .C1(G234), .C2(G237), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT14), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n188), .A2(G122), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n428), .B(new_n430), .C1(new_n193), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n188), .A2(KEYINPUT69), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G116), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n437), .A3(G107), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n299), .B(new_n430), .C1(new_n193), .C2(new_n431), .ZN(new_n439));
  XOR2_X1   g253(.A(G128), .B(G143), .Z(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G134), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n440), .A2(G134), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n438), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G107), .B1(new_n436), .B2(new_n429), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n439), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT13), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n202), .A3(G128), .ZN(new_n447));
  OAI211_X1 g261(.A(G134), .B(new_n447), .C1(new_n440), .C2(new_n446), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT94), .B1(new_n440), .B2(G134), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n440), .A2(KEYINPUT94), .A3(G134), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT9), .B(G234), .ZN(new_n453));
  INV_X1    g267(.A(G217), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n453), .A2(new_n454), .A3(G953), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n443), .A2(new_n451), .A3(new_n455), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n452), .A2(KEYINPUT95), .A3(new_n456), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n187), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G478), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT15), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n460), .A2(new_n187), .A3(new_n461), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n417), .A2(new_n427), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G221), .B1(new_n453), .B2(G902), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G469), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n187), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n312), .A2(new_n242), .A3(new_n314), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n319), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n475));
  INV_X1    g289(.A(new_n237), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n213), .A2(new_n311), .A3(new_n317), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT10), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n213), .B1(new_n311), .B2(new_n317), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n476), .B1(new_n481), .B2(KEYINPUT81), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT12), .B1(new_n237), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n318), .A2(new_n333), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n477), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n482), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n485), .B1(new_n482), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G140), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n336), .A2(G227), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n480), .A2(new_n494), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n237), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n491), .A2(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n473), .B1(new_n499), .B2(G469), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n480), .A2(new_n494), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n482), .A2(new_n485), .A3(new_n488), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n484), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n494), .B1(new_n498), .B2(new_n480), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n472), .B(new_n187), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(KEYINPUT83), .B(new_n471), .C1(new_n500), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n496), .A2(new_n498), .ZN(new_n510));
  INV_X1    g324(.A(new_n497), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n504), .A2(new_n502), .B1(new_n511), .B2(new_n476), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(G469), .C1(new_n512), .C2(new_n494), .ZN(new_n513));
  INV_X1    g327(.A(new_n473), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n509), .B1(new_n515), .B2(new_n470), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n360), .B(new_n469), .C1(new_n508), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n454), .B1(G234), .B2(new_n187), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT74), .B1(new_n194), .B2(G128), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n520), .A2(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n194), .A2(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(KEYINPUT23), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G110), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT73), .B1(new_n194), .B2(G128), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n198), .A3(G119), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n528), .A2(new_n530), .B1(new_n194), .B2(G128), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT24), .B(G110), .Z(new_n532));
  OAI21_X1  g346(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR3_X1    g347(.A1(new_n531), .A2(new_n527), .A3(new_n532), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n526), .A2(new_n537), .A3(new_n533), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n363), .A2(new_n200), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n536), .A2(new_n365), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n378), .A2(new_n365), .B1(new_n531), .B2(new_n532), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n525), .B2(new_n524), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n336), .A2(G221), .A3(G234), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT22), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(G137), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n542), .A3(new_n546), .ZN(new_n549));
  XOR2_X1   g363(.A(KEYINPUT77), .B(KEYINPUT25), .Z(new_n550));
  NAND4_X1  g364(.A1(new_n548), .A2(new_n187), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n540), .A2(new_n542), .A3(new_n546), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n546), .B1(new_n540), .B2(new_n542), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n519), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT78), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n548), .A2(new_n558), .A3(new_n549), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n519), .A2(G902), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n295), .A2(new_n518), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  INV_X1    g379(.A(new_n360), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n460), .A2(new_n567), .A3(new_n461), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n457), .A2(KEYINPUT33), .A3(new_n459), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n568), .A2(new_n569), .A3(G478), .A4(new_n187), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n462), .A2(new_n463), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n417), .A2(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n566), .A2(new_n427), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G472), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n289), .B2(new_n187), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n269), .B2(new_n289), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n508), .A2(new_n516), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n574), .A2(new_n577), .A3(new_n563), .A4(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT34), .B(G104), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT97), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(G6));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n416), .B1(new_n408), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n408), .A2(new_n584), .A3(new_n410), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n426), .B(KEYINPUT99), .Z(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n586), .A2(new_n468), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n590), .A2(KEYINPUT100), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(KEYINPUT100), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n360), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n579), .A2(new_n563), .A3(new_n577), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT35), .B(G107), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G9));
  NOR2_X1   g411(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n543), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n560), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n556), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n518), .A2(new_n577), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT37), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n525), .ZN(G12));
  INV_X1    g418(.A(new_n508), .ZN(new_n605));
  INV_X1    g419(.A(new_n516), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n566), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n587), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n585), .ZN(new_n609));
  INV_X1    g423(.A(G900), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n421), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n425), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n609), .A2(new_n468), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n295), .A2(new_n607), .A3(new_n601), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT101), .B(G128), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G30));
  INV_X1    g430(.A(new_n277), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n258), .A2(new_n259), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n281), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n619), .B2(G902), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n291), .B2(new_n294), .ZN(new_n621));
  INV_X1    g435(.A(new_n601), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n415), .B1(new_n408), .B2(new_n410), .ZN(new_n623));
  INV_X1    g437(.A(new_n297), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n468), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n358), .A2(new_n359), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT38), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n621), .A2(new_n622), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n629), .A2(KEYINPUT102), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n612), .B(KEYINPUT39), .Z(new_n631));
  NOR2_X1   g445(.A1(new_n578), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(KEYINPUT102), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G143), .ZN(G45));
  AOI22_X1  g450(.A1(new_n411), .A2(new_n416), .B1(new_n571), .B2(new_n570), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n637), .A2(KEYINPUT103), .A3(new_n612), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT103), .B1(new_n637), .B2(new_n612), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n295), .A2(new_n607), .A3(new_n601), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G146), .ZN(G48));
  OR2_X1    g456(.A1(new_n505), .A2(new_n506), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n187), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G469), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n470), .A3(new_n507), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT104), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n645), .A2(new_n648), .A3(new_n470), .A4(new_n507), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n295), .A2(new_n563), .A3(new_n574), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  NAND2_X1  g467(.A1(new_n295), .A2(new_n563), .ZN(new_n654));
  INV_X1    g468(.A(new_n650), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n593), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT105), .B(G116), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G18));
  NOR2_X1   g472(.A1(new_n646), .A2(new_n566), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n295), .A2(new_n469), .A3(new_n601), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G119), .ZN(G21));
  AOI21_X1  g475(.A(new_n588), .B1(new_n647), .B2(new_n649), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n626), .A2(new_n627), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n664));
  INV_X1    g478(.A(new_n269), .ZN(new_n665));
  AOI22_X1  g479(.A1(KEYINPUT31), .A2(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n666), .A2(new_n667), .B1(new_n272), .B2(new_n617), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n278), .A2(new_n282), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT106), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n576), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n664), .B1(new_n672), .B2(new_n563), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n576), .A2(new_n671), .A3(new_n562), .A4(KEYINPUT107), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n662), .B(new_n663), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  NOR3_X1   g490(.A1(new_n622), .A2(new_n576), .A3(new_n671), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n640), .A2(new_n659), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT108), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n331), .ZN(G27));
  NAND2_X1  g494(.A1(new_n515), .A2(KEYINPUT109), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n500), .A2(new_n682), .A3(new_n507), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n471), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n627), .A2(new_n297), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n295), .A2(new_n563), .A3(new_n686), .A4(new_n640), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n292), .A2(new_n293), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(new_n268), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n562), .B1(new_n691), .B2(new_n285), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n640), .A4(new_n686), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G131), .ZN(G33));
  AND4_X1   g509(.A1(new_n563), .A2(new_n295), .A3(new_n613), .A4(new_n686), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n216), .ZN(G36));
  NAND2_X1  g511(.A1(new_n623), .A2(new_n572), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT43), .ZN(new_n699));
  OR3_X1    g513(.A1(new_n577), .A2(new_n699), .A3(new_n622), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n297), .B(new_n627), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n499), .B(KEYINPUT45), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT46), .B1(new_n704), .B2(new_n514), .ZN(new_n705));
  INV_X1    g519(.A(new_n507), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n704), .A2(KEYINPUT46), .A3(new_n514), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n471), .A3(new_n631), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n702), .B(new_n710), .C1(new_n701), .C2(new_n700), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G137), .ZN(G39));
  OAI22_X1  g526(.A1(new_n709), .A2(new_n471), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n709), .B2(new_n471), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n690), .A2(new_n286), .A3(new_n285), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n287), .A2(new_n290), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n268), .A2(new_n640), .A3(new_n722), .A4(new_n685), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n718), .A2(new_n719), .A3(new_n562), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G140), .ZN(G42));
  NAND2_X1  g539(.A1(new_n645), .A2(new_n507), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n563), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n729), .A2(new_n471), .A3(new_n297), .A4(new_n698), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n730), .A2(new_n731), .B1(new_n728), .B2(new_n727), .ZN(new_n733));
  INV_X1    g547(.A(new_n621), .ZN(new_n734));
  INV_X1    g548(.A(new_n628), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n732), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n726), .A2(new_n470), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n718), .B2(new_n719), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n673), .A2(new_n674), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n699), .A2(new_n425), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n685), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT51), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n727), .A2(new_n685), .A3(new_n470), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT118), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n740), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n677), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n563), .A3(new_n424), .A4(new_n734), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n749), .A2(new_n417), .A3(new_n572), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n741), .A2(new_n646), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n628), .A2(new_n624), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(KEYINPUT50), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT50), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n748), .B(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(G952), .B(new_n336), .C1(new_n744), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n718), .A2(new_n719), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n737), .B(KEYINPUT117), .Z(new_n759));
  OAI211_X1 g573(.A(new_n685), .B(new_n742), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n753), .A2(new_n754), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n748), .A4(new_n750), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n756), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n623), .A2(new_n468), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n573), .A2(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n765), .A2(new_n360), .A3(new_n589), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n579), .A3(new_n577), .A4(new_n563), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n564), .A2(new_n602), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n564), .A2(new_n602), .A3(new_n767), .A4(KEYINPUT112), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n656), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n696), .B1(new_n689), .B2(new_n693), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n675), .A2(new_n651), .A3(new_n660), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n772), .A2(new_n773), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n686), .A2(new_n640), .A3(new_n677), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n622), .B1(new_n722), .B2(new_n268), .ZN(new_n780));
  INV_X1    g594(.A(new_n468), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n685), .A2(new_n781), .A3(new_n609), .A4(new_n612), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n578), .B1(new_n782), .B2(KEYINPUT113), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n780), .B(new_n783), .C1(KEYINPUT113), .C2(new_n782), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT114), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n777), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n684), .A2(new_n663), .A3(new_n612), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n621), .A2(new_n787), .A3(new_n622), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n614), .A2(new_n641), .A3(new_n788), .A4(new_n678), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n780), .B(new_n607), .C1(new_n613), .C2(new_n640), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n678), .A4(new_n788), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT116), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n790), .B2(new_n793), .ZN(new_n800));
  INV_X1    g614(.A(new_n797), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n786), .A2(KEYINPUT53), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n656), .B(new_n775), .C1(new_n770), .C2(new_n771), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n784), .B(KEYINPUT114), .Z(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n778), .A4(new_n774), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n790), .A2(new_n793), .A3(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n796), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n804), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n803), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n807), .A2(new_n809), .A3(new_n804), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n786), .A2(new_n802), .A3(new_n798), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n813), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n763), .B(new_n812), .C1(new_n815), .C2(new_n811), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n749), .A2(new_n573), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n741), .A2(new_n566), .A3(new_n646), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n747), .A2(new_n692), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT48), .Z(new_n820));
  NOR4_X1   g634(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(G952), .A2(G953), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n736), .B1(new_n821), .B2(new_n822), .ZN(G75));
  XOR2_X1   g637(.A(new_n338), .B(KEYINPUT120), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n330), .A2(new_n340), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT119), .Z(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT55), .Z(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n187), .B1(new_n803), .B2(new_n810), .ZN(new_n829));
  AOI211_X1 g643(.A(KEYINPUT56), .B(new_n828), .C1(new_n829), .C2(G210), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n803), .A2(new_n810), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(G210), .A3(G902), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n827), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n824), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n336), .A2(G952), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(G210), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n838), .B(new_n187), .C1(new_n803), .C2(new_n810), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n828), .B1(new_n839), .B2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n833), .A3(new_n827), .ZN(new_n841));
  INV_X1    g655(.A(new_n824), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n835), .A2(new_n837), .A3(new_n843), .ZN(G51));
  NAND2_X1  g658(.A1(new_n514), .A2(KEYINPUT57), .ZN(new_n845));
  INV_X1    g659(.A(new_n812), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n811), .B1(new_n803), .B2(new_n810), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n514), .A2(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n643), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n829), .A2(G469), .A3(new_n703), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n836), .B1(new_n850), .B2(new_n851), .ZN(G54));
  NAND3_X1  g666(.A1(new_n829), .A2(KEYINPUT58), .A3(G475), .ZN(new_n853));
  INV_X1    g667(.A(new_n405), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n856), .A3(new_n836), .ZN(G60));
  NAND2_X1  g671(.A1(new_n568), .A2(new_n569), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n812), .B1(new_n815), .B2(new_n811), .ZN(new_n860));
  NAND2_X1  g674(.A1(G478), .A2(G902), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT59), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n859), .B(new_n862), .C1(new_n846), .C2(new_n847), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n863), .A2(new_n865), .A3(new_n836), .ZN(G63));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n867));
  NAND2_X1  g681(.A1(G217), .A2(G902), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT60), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n803), .B2(new_n810), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n557), .A2(new_n559), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT121), .B1(new_n872), .B2(new_n837), .ZN(new_n873));
  OAI211_X1 g687(.A(KEYINPUT121), .B(new_n837), .C1(new_n870), .C2(new_n871), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n599), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n867), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n870), .A2(new_n871), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n878), .A2(KEYINPUT122), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n867), .B1(new_n878), .B2(KEYINPUT122), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n837), .A4(new_n875), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(G66));
  AOI21_X1  g696(.A(new_n336), .B1(new_n419), .B2(G224), .ZN(new_n883));
  INV_X1    g697(.A(new_n805), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n336), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n826), .B1(G898), .B2(new_n336), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT123), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n885), .B(new_n887), .ZN(G69));
  NAND3_X1  g702(.A1(new_n710), .A2(new_n663), .A3(new_n692), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n889), .A2(new_n774), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n791), .A2(new_n678), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n711), .A3(new_n724), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n336), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n245), .A2(new_n246), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n398), .A2(new_n399), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n893), .B(new_n897), .C1(G900), .C2(new_n336), .ZN(new_n898));
  INV_X1    g712(.A(new_n654), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n632), .A3(new_n685), .A4(new_n765), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n724), .A2(new_n711), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n635), .B(new_n891), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n635), .A2(new_n891), .A3(new_n902), .A4(new_n903), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n336), .A3(new_n896), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n336), .B1(G227), .B2(G900), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT125), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n898), .A2(new_n908), .B1(KEYINPUT126), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(KEYINPUT126), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G72));
  NAND2_X1  g727(.A1(G472), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT63), .Z(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n907), .B2(new_n884), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n251), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n256), .C1(new_n917), .C2(new_n916), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n892), .B2(new_n884), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n281), .A3(new_n251), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n837), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n915), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n257), .A2(new_n617), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n815), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G57));
endmodule


