

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n731), .ZN(n695) );
  AND2_X1 U552 ( .A1(n950), .A2(n808), .ZN(n517) );
  AND2_X1 U553 ( .A1(n695), .A2(G1996), .ZN(n681) );
  INV_X1 U554 ( .A(KEYINPUT97), .ZN(n693) );
  XNOR2_X1 U555 ( .A(n694), .B(n693), .ZN(n701) );
  NOR2_X1 U556 ( .A1(n794), .A2(n517), .ZN(n795) );
  NOR2_X1 U557 ( .A1(G2105), .A2(n537), .ZN(n870) );
  NOR2_X1 U558 ( .A1(G651), .A2(n646), .ZN(n641) );
  XNOR2_X1 U559 ( .A(n549), .B(KEYINPUT86), .ZN(G164) );
  INV_X1 U560 ( .A(G651), .ZN(n523) );
  NOR2_X1 U561 ( .A1(G543), .A2(n523), .ZN(n518) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n518), .Z(n645) );
  NAND2_X1 U563 ( .A1(G63), .A2(n645), .ZN(n520) );
  XOR2_X1 U564 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  NAND2_X1 U565 ( .A1(G51), .A2(n641), .ZN(n519) );
  NAND2_X1 U566 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U567 ( .A(KEYINPUT6), .B(n521), .ZN(n529) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n635) );
  NAND2_X1 U569 ( .A1(n635), .A2(G89), .ZN(n522) );
  XNOR2_X1 U570 ( .A(n522), .B(KEYINPUT4), .ZN(n526) );
  OR2_X1 U571 ( .A1(n523), .A2(n646), .ZN(n524) );
  XNOR2_X1 U572 ( .A(KEYINPUT67), .B(n524), .ZN(n632) );
  NAND2_X1 U573 ( .A1(G76), .A2(n632), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U575 ( .A(n527), .B(KEYINPUT5), .Z(n528) );
  NOR2_X1 U576 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U577 ( .A(KEYINPUT7), .B(n530), .Z(n532) );
  XOR2_X1 U578 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n531) );
  XNOR2_X1 U579 ( .A(n532), .B(n531), .ZN(G168) );
  XOR2_X1 U580 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT65), .ZN(n867) );
  NAND2_X1 U583 ( .A1(n867), .A2(G113), .ZN(n536) );
  INV_X1 U584 ( .A(G2104), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G101), .A2(n870), .ZN(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n534), .Z(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n542) );
  AND2_X1 U588 ( .A1(n537), .A2(G2105), .ZN(n866) );
  NAND2_X1 U589 ( .A1(G125), .A2(n866), .ZN(n540) );
  NOR2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n538), .Z(n871) );
  NAND2_X1 U592 ( .A1(G137), .A2(n871), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X2 U594 ( .A1(n542), .A2(n541), .ZN(G160) );
  NAND2_X1 U595 ( .A1(G102), .A2(n870), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G138), .A2(n871), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U598 ( .A1(G126), .A2(n866), .ZN(n546) );
  NAND2_X1 U599 ( .A1(G114), .A2(n867), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G64), .A2(n645), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G52), .A2(n641), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U605 ( .A1(n632), .A2(G77), .ZN(n553) );
  NAND2_X1 U606 ( .A1(n635), .A2(G90), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U609 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  XOR2_X1 U613 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n558) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(G223) );
  INV_X1 U616 ( .A(G223), .ZN(n813) );
  NAND2_X1 U617 ( .A1(n813), .A2(G567), .ZN(n559) );
  XOR2_X1 U618 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U619 ( .A1(G56), .A2(n645), .ZN(n560) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(n560), .Z(n567) );
  NAND2_X1 U621 ( .A1(G81), .A2(n635), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n561), .B(KEYINPUT70), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G68), .A2(n632), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n565), .Z(n566) );
  NOR2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n641), .A2(G43), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n929) );
  XNOR2_X1 U630 ( .A(G860), .B(KEYINPUT71), .ZN(n589) );
  OR2_X1 U631 ( .A1(n929), .A2(n589), .ZN(G153) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  INV_X1 U633 ( .A(G868), .ZN(n659) );
  NAND2_X1 U634 ( .A1(G92), .A2(n635), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G66), .A2(n645), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G79), .A2(n632), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G54), .A2(n641), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT15), .B(n576), .Z(n945) );
  AND2_X1 U642 ( .A1(n659), .A2(n945), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n659), .A2(G301), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT72), .B(n579), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G65), .A2(n645), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G53), .A2(n641), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G91), .A2(n635), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G78), .A2(n632), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n946) );
  INV_X1 U653 ( .A(n946), .ZN(G299) );
  NAND2_X1 U654 ( .A1(G299), .A2(n659), .ZN(n587) );
  NAND2_X1 U655 ( .A1(G868), .A2(G286), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT75), .B(n588), .Z(G297) );
  NAND2_X1 U658 ( .A1(n589), .A2(G559), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n590), .A2(n945), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U661 ( .A1(G868), .A2(n929), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G868), .A2(n945), .ZN(n592) );
  NOR2_X1 U663 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U665 ( .A1(G123), .A2(n866), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT76), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(KEYINPUT18), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G111), .A2(n867), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G99), .A2(n870), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G135), .A2(n871), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT77), .B(n603), .Z(n1000) );
  XNOR2_X1 U675 ( .A(n1000), .B(G2096), .ZN(n605) );
  INV_X1 U676 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U678 ( .A1(G559), .A2(n945), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(n929), .ZN(n656) );
  NOR2_X1 U680 ( .A1(n656), .A2(G860), .ZN(n614) );
  NAND2_X1 U681 ( .A1(G55), .A2(n641), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT78), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n645), .A2(G67), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G93), .A2(n635), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G80), .A2(n632), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n658) );
  XOR2_X1 U689 ( .A(n614), .B(n658), .Z(G145) );
  NAND2_X1 U690 ( .A1(G75), .A2(n632), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT82), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n645), .A2(G62), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G50), .A2(n641), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G88), .A2(n635), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT81), .B(n619), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(G303) );
  INV_X1 U700 ( .A(G303), .ZN(G166) );
  NAND2_X1 U701 ( .A1(G86), .A2(n635), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G48), .A2(n641), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G73), .A2(n632), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n626), .B(KEYINPUT2), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n627), .B(KEYINPUT79), .ZN(n628) );
  NOR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n645), .A2(G61), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G72), .A2(n632), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G60), .A2(n645), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n635), .A2(G85), .ZN(n636) );
  XOR2_X1 U714 ( .A(KEYINPUT66), .B(n636), .Z(n637) );
  NOR2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(G47), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(G290) );
  NAND2_X1 U718 ( .A1(G49), .A2(n641), .ZN(n643) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(G288) );
  XOR2_X1 U724 ( .A(n658), .B(KEYINPUT19), .Z(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(KEYINPUT83), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n946), .B(G305), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n650), .B(G290), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U730 ( .A(G166), .B(n654), .ZN(n885) );
  XOR2_X1 U731 ( .A(n885), .B(KEYINPUT84), .Z(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U742 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U745 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U746 ( .A1(G96), .A2(n668), .ZN(n818) );
  NAND2_X1 U747 ( .A1(n818), .A2(G2106), .ZN(n672) );
  NAND2_X1 U748 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U749 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G108), .A2(n670), .ZN(n819) );
  NAND2_X1 U751 ( .A1(n819), .A2(G567), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n672), .A2(n671), .ZN(n839) );
  NAND2_X1 U753 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U754 ( .A1(n839), .A2(n673), .ZN(n816) );
  NAND2_X1 U755 ( .A1(n816), .A2(G36), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT85), .B(n674), .Z(G176) );
  NAND2_X1 U757 ( .A1(G160), .A2(G40), .ZN(n779) );
  INV_X1 U758 ( .A(n779), .ZN(n675) );
  NOR2_X1 U759 ( .A1(G1384), .A2(G164), .ZN(n780) );
  NAND2_X2 U760 ( .A1(n675), .A2(n780), .ZN(n731) );
  NAND2_X1 U761 ( .A1(G8), .A2(n731), .ZN(n754) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n676) );
  XOR2_X1 U763 ( .A(n676), .B(KEYINPUT24), .Z(n677) );
  NOR2_X1 U764 ( .A1(n754), .A2(n677), .ZN(n759) );
  INV_X1 U765 ( .A(G1961), .ZN(n956) );
  NAND2_X1 U766 ( .A1(n731), .A2(n956), .ZN(n679) );
  XNOR2_X1 U767 ( .A(KEYINPUT25), .B(G2078), .ZN(n907) );
  NAND2_X1 U768 ( .A1(n695), .A2(n907), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n715) );
  NAND2_X1 U770 ( .A1(n715), .A2(G171), .ZN(n709) );
  XOR2_X1 U771 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n680) );
  XNOR2_X1 U772 ( .A(n681), .B(n680), .ZN(n684) );
  AND2_X1 U773 ( .A1(n731), .A2(G1341), .ZN(n682) );
  NOR2_X1 U774 ( .A1(n682), .A2(n929), .ZN(n683) );
  AND2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n685) );
  OR2_X1 U776 ( .A1(n945), .A2(n685), .ZN(n692) );
  NAND2_X1 U777 ( .A1(n685), .A2(n945), .ZN(n690) );
  INV_X1 U778 ( .A(G2067), .ZN(n909) );
  NOR2_X1 U779 ( .A1(n731), .A2(n909), .ZN(n686) );
  XOR2_X1 U780 ( .A(n686), .B(KEYINPUT96), .Z(n688) );
  NAND2_X1 U781 ( .A1(n731), .A2(G1348), .ZN(n687) );
  NAND2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n731), .A2(G1956), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n695), .A2(G2072), .ZN(n696) );
  XOR2_X1 U787 ( .A(KEYINPUT27), .B(n696), .Z(n697) );
  NAND2_X1 U788 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT95), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n702), .A2(n946), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U792 ( .A1(n702), .A2(n946), .ZN(n703) );
  XOR2_X1 U793 ( .A(n703), .B(KEYINPUT28), .Z(n704) );
  NAND2_X1 U794 ( .A1(n705), .A2(n704), .ZN(n707) );
  XOR2_X1 U795 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n706) );
  XNOR2_X1 U796 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n720) );
  NOR2_X1 U798 ( .A1(n754), .A2(G1966), .ZN(n710) );
  XNOR2_X1 U799 ( .A(n710), .B(KEYINPUT94), .ZN(n721) );
  NOR2_X1 U800 ( .A1(n731), .A2(G2084), .ZN(n711) );
  XNOR2_X1 U801 ( .A(n711), .B(KEYINPUT93), .ZN(n722) );
  NAND2_X1 U802 ( .A1(G8), .A2(n722), .ZN(n712) );
  NOR2_X1 U803 ( .A1(n721), .A2(n712), .ZN(n713) );
  XOR2_X1 U804 ( .A(KEYINPUT30), .B(n713), .Z(n714) );
  NOR2_X1 U805 ( .A1(G168), .A2(n714), .ZN(n717) );
  NOR2_X1 U806 ( .A1(G171), .A2(n715), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U808 ( .A(KEYINPUT31), .B(n718), .Z(n719) );
  NAND2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n729) );
  INV_X1 U810 ( .A(n729), .ZN(n727) );
  INV_X1 U811 ( .A(n721), .ZN(n725) );
  INV_X1 U812 ( .A(n722), .ZN(n723) );
  NAND2_X1 U813 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U815 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U816 ( .A(KEYINPUT99), .B(n728), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n729), .A2(G286), .ZN(n736) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n754), .ZN(n730) );
  XNOR2_X1 U819 ( .A(n730), .B(KEYINPUT100), .ZN(n733) );
  NOR2_X1 U820 ( .A1(n731), .A2(G2090), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n734), .A2(G303), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U825 ( .A(n738), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n753) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n746) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U829 ( .A1(n746), .A2(n741), .ZN(n933) );
  XOR2_X1 U830 ( .A(n933), .B(KEYINPUT101), .Z(n742) );
  NAND2_X1 U831 ( .A1(n753), .A2(n742), .ZN(n743) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NAND2_X1 U833 ( .A1(n743), .A2(n932), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n754), .A2(n744), .ZN(n745) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n745), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n746), .A2(KEYINPUT33), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n747), .A2(n754), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n941) );
  NAND2_X1 U840 ( .A1(n750), .A2(n941), .ZN(n757) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U842 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  INV_X1 U847 ( .A(n760), .ZN(n796) );
  NAND2_X1 U848 ( .A1(G141), .A2(n871), .ZN(n761) );
  XNOR2_X1 U849 ( .A(n761), .B(KEYINPUT90), .ZN(n768) );
  NAND2_X1 U850 ( .A1(G129), .A2(n866), .ZN(n763) );
  NAND2_X1 U851 ( .A1(G117), .A2(n867), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n870), .A2(G105), .ZN(n764) );
  XOR2_X1 U854 ( .A(KEYINPUT38), .B(n764), .Z(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n877) );
  NAND2_X1 U857 ( .A1(G1996), .A2(n877), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n769), .B(KEYINPUT91), .ZN(n778) );
  NAND2_X1 U859 ( .A1(G119), .A2(n866), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G107), .A2(n867), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G95), .A2(n870), .ZN(n772) );
  XNOR2_X1 U863 ( .A(KEYINPUT89), .B(n772), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n871), .A2(G131), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n863) );
  AND2_X1 U867 ( .A1(G1991), .A2(n863), .ZN(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n991) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n808) );
  XOR2_X1 U870 ( .A(n808), .B(KEYINPUT92), .Z(n781) );
  NOR2_X1 U871 ( .A1(n991), .A2(n781), .ZN(n800) );
  INV_X1 U872 ( .A(n800), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G104), .A2(n870), .ZN(n783) );
  NAND2_X1 U874 ( .A1(G140), .A2(n871), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n784) );
  XNOR2_X1 U877 ( .A(n785), .B(n784), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n866), .A2(G128), .ZN(n786) );
  XNOR2_X1 U879 ( .A(n786), .B(KEYINPUT88), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G116), .A2(n867), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U882 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U884 ( .A(KEYINPUT36), .B(n792), .ZN(n850) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NOR2_X1 U886 ( .A1(n850), .A2(n805), .ZN(n993) );
  NAND2_X1 U887 ( .A1(n808), .A2(n993), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n793), .A2(n803), .ZN(n794) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n950) );
  NAND2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n811) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n877), .ZN(n987) );
  NOR2_X1 U892 ( .A1(n863), .A2(G1991), .ZN(n797) );
  XNOR2_X1 U893 ( .A(n797), .B(KEYINPUT102), .ZN(n999) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n999), .A2(n798), .ZN(n799) );
  NOR2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U897 ( .A1(n987), .A2(n801), .ZN(n802) );
  XNOR2_X1 U898 ( .A(n802), .B(KEYINPUT39), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n850), .A2(n805), .ZN(n989) );
  NAND2_X1 U901 ( .A1(n806), .A2(n989), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U903 ( .A(KEYINPUT103), .B(n809), .Z(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U905 ( .A(KEYINPUT40), .B(n812), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n815) );
  XNOR2_X1 U910 ( .A(KEYINPUT106), .B(n815), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(G188) );
  INV_X1 U913 ( .A(G120), .ZN(G236) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  XOR2_X1 U918 ( .A(KEYINPUT107), .B(G2090), .Z(n821) );
  XNOR2_X1 U919 ( .A(G2067), .B(G2084), .ZN(n820) );
  XNOR2_X1 U920 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U921 ( .A(n822), .B(G2100), .Z(n824) );
  XNOR2_X1 U922 ( .A(G2078), .B(G2072), .ZN(n823) );
  XNOR2_X1 U923 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U924 ( .A(G2096), .B(G2678), .Z(n826) );
  XNOR2_X1 U925 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U927 ( .A(n828), .B(n827), .Z(G227) );
  XNOR2_X1 U928 ( .A(G1981), .B(KEYINPUT108), .ZN(n838) );
  XOR2_X1 U929 ( .A(G1976), .B(G1956), .Z(n830) );
  XNOR2_X1 U930 ( .A(G1966), .B(G1961), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U932 ( .A(G1986), .B(G1971), .Z(n832) );
  XNOR2_X1 U933 ( .A(G1991), .B(G1996), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U935 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U936 ( .A(G2474), .B(KEYINPUT41), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G229) );
  INV_X1 U939 ( .A(n839), .ZN(G319) );
  NAND2_X1 U940 ( .A1(n866), .A2(G124), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n840), .B(KEYINPUT44), .ZN(n842) );
  NAND2_X1 U942 ( .A1(G112), .A2(n867), .ZN(n841) );
  NAND2_X1 U943 ( .A1(n842), .A2(n841), .ZN(n846) );
  NAND2_X1 U944 ( .A1(G100), .A2(n870), .ZN(n844) );
  NAND2_X1 U945 ( .A1(G136), .A2(n871), .ZN(n843) );
  NAND2_X1 U946 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U947 ( .A1(n846), .A2(n845), .ZN(G162) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(KEYINPUT112), .ZN(n848) );
  XNOR2_X1 U949 ( .A(G164), .B(G160), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U951 ( .A(KEYINPUT46), .B(n849), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n850), .B(KEYINPUT48), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n853), .B(G162), .Z(n865) );
  NAND2_X1 U955 ( .A1(G103), .A2(n870), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G139), .A2(n871), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n862) );
  NAND2_X1 U958 ( .A1(n866), .A2(G127), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n856), .B(KEYINPUT110), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G115), .A2(n867), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U962 ( .A(KEYINPUT47), .B(n859), .ZN(n860) );
  XNOR2_X1 U963 ( .A(KEYINPUT111), .B(n860), .ZN(n861) );
  NOR2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n994) );
  XOR2_X1 U965 ( .A(n863), .B(n994), .Z(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n881) );
  NAND2_X1 U967 ( .A1(G130), .A2(n866), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G118), .A2(n867), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G106), .A2(n870), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G142), .A2(n871), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U973 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(n1000), .B(n879), .Z(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U978 ( .A1(G37), .A2(n882), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n929), .B(KEYINPUT113), .ZN(n884) );
  XNOR2_X1 U980 ( .A(G171), .B(n945), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n887) );
  XOR2_X1 U982 ( .A(G286), .B(n885), .Z(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U984 ( .A1(G37), .A2(n888), .ZN(G397) );
  XNOR2_X1 U985 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n890) );
  NOR2_X1 U986 ( .A1(G227), .A2(G229), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n903) );
  XNOR2_X1 U988 ( .A(G2446), .B(KEYINPUT104), .ZN(n900) );
  XOR2_X1 U989 ( .A(KEYINPUT105), .B(G2427), .Z(n892) );
  XNOR2_X1 U990 ( .A(G2435), .B(G2438), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U992 ( .A(G2454), .B(G2430), .Z(n894) );
  XNOR2_X1 U993 ( .A(G1341), .B(G1348), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2451), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n901), .A2(G14), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n906), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  INV_X1 U1006 ( .A(n906), .ZN(G401) );
  XNOR2_X1 U1007 ( .A(G27), .B(n907), .ZN(n919) );
  XNOR2_X1 U1008 ( .A(G25), .B(G1991), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n908), .B(KEYINPUT119), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(G26), .B(n909), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n910), .A2(G28), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(G33), .B(G2072), .ZN(n911) );
  NOR2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT120), .B(G1996), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(G32), .B(n915), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n920), .B(KEYINPUT53), .ZN(n923) );
  XOR2_X1 U1020 ( .A(G2084), .B(KEYINPUT54), .Z(n921) );
  XNOR2_X1 U1021 ( .A(G34), .B(n921), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT118), .B(G2090), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G35), .B(n924), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1026 ( .A(KEYINPUT55), .B(n927), .Z(n928) );
  NOR2_X1 U1027 ( .A1(G29), .A2(n928), .ZN(n984) );
  XNOR2_X1 U1028 ( .A(G16), .B(KEYINPUT56), .ZN(n954) );
  XNOR2_X1 U1029 ( .A(G301), .B(G1961), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n929), .B(G1341), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n938) );
  AND2_X1 U1032 ( .A1(G303), .A2(G1971), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n936), .B(KEYINPUT122), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n944) );
  XOR2_X1 U1037 ( .A(G1966), .B(KEYINPUT121), .Z(n939) );
  XNOR2_X1 U1038 ( .A(G168), .B(n939), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1040 ( .A(KEYINPUT57), .B(n942), .Z(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1042 ( .A(n945), .B(G1348), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n946), .B(G1956), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n955), .B(KEYINPUT123), .ZN(n981) );
  XOR2_X1 U1049 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n977) );
  XOR2_X1 U1050 ( .A(G1966), .B(G21), .Z(n958) );
  XNOR2_X1 U1051 ( .A(n956), .B(G5), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n975) );
  XOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .Z(n966) );
  XNOR2_X1 U1061 ( .A(G4), .B(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(G20), .B(G1956), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1068 ( .A(KEYINPUT60), .B(n973), .Z(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(KEYINPUT124), .B(n978), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n979), .A2(G16), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n982), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n985), .B(KEYINPUT126), .ZN(n1016) );
  XOR2_X1 U1077 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT51), .B(n988), .Z(n990) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n1010) );
  INV_X1 U1081 ( .A(n991), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n1008) );
  XOR2_X1 U1083 ( .A(G2072), .B(n994), .Z(n996) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1086 ( .A(KEYINPUT50), .B(n997), .Z(n1006) );
  XNOR2_X1 U1087 ( .A(G160), .B(G2084), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT115), .ZN(n1003) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT116), .B(n1001), .Z(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(KEYINPUT117), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1011), .ZN(n1013) );
  INV_X1 U1097 ( .A(KEYINPUT55), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

