//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  OR3_X1    g0016(.A1(new_n215), .A2(new_n209), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n216), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(new_n252), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n255), .A2(KEYINPUT66), .A3(new_n248), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n254), .A2(new_n256), .B1(G1), .B2(new_n209), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n250), .B1(new_n257), .B2(new_n247), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT72), .B1(new_n202), .B2(new_n203), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT72), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G58), .A3(G68), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n259), .B(new_n261), .C1(G58), .C2(G68), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n262), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT70), .B(KEYINPUT3), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n209), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n268), .A2(new_n270), .B1(new_n274), .B2(new_n269), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n264), .B1(new_n275), .B2(new_n203), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT16), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n255), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G33), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT71), .B1(new_n271), .B2(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT71), .A4(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n209), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n284), .A2(new_n269), .A3(new_n209), .A4(new_n285), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G68), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT16), .B(new_n264), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n258), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G226), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G1698), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G223), .B2(G1698), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n284), .B2(new_n285), .ZN(new_n296));
  INV_X1    g0096(.A(G87), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n271), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n292), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n292), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  OAI211_X1 g0103(.A(G1), .B(G13), .C1(new_n271), .C2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n304), .A2(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n302), .B1(G232), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n299), .A2(G190), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n299), .B2(new_n306), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n291), .A2(new_n310), .A3(KEYINPUT74), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT17), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n278), .A2(new_n290), .ZN(new_n313));
  INV_X1    g0113(.A(new_n258), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n299), .A2(new_n306), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n317), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT18), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT18), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n317), .A2(new_n325), .A3(new_n318), .A4(new_n322), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n312), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G1698), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n273), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(G223), .B1(G77), .B2(new_n273), .ZN(new_n331));
  INV_X1    g0131(.A(G222), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n272), .A2(new_n266), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n329), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n292), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n302), .B1(G226), .B2(new_n305), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n257), .A2(new_n201), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n271), .A2(G20), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n247), .A2(new_n342), .B1(G150), .B2(new_n263), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n204), .A2(G20), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n255), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT65), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(new_n346), .B1(new_n201), .B2(new_n249), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n336), .A2(new_n321), .A3(new_n337), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n340), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT68), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n338), .B2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n336), .A2(KEYINPUT68), .A3(G190), .A4(new_n337), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(new_n356), .B1(G200), .B2(new_n338), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n349), .A2(KEYINPUT67), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT67), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n341), .A2(new_n347), .A3(new_n348), .A4(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(KEYINPUT9), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT9), .B1(new_n358), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT10), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n363), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n361), .A4(new_n357), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n352), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n342), .A2(G77), .ZN(new_n369));
  INV_X1    g0169(.A(new_n263), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n369), .B1(new_n209), .B2(G68), .C1(new_n201), .C2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n249), .A2(new_n203), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n253), .B(G68), .C1(G1), .C2(new_n209), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT11), .B1(new_n371), .B2(new_n252), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT14), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G97), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n334), .B2(new_n293), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n273), .A2(new_n231), .A3(new_n329), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n292), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n302), .B1(G238), .B2(new_n305), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n379), .B(G169), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n383), .A2(new_n385), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(G179), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n386), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n379), .B1(new_n394), .B2(G169), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n378), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n387), .A2(new_n388), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n378), .B1(new_n397), .B2(G190), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT69), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(G200), .C1(new_n387), .C2(new_n388), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n394), .B2(G200), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n247), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n297), .A2(KEYINPUT15), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT15), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G87), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n342), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n255), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n253), .ZN(new_n411));
  OAI21_X1  g0211(.A(G77), .B1(new_n209), .B2(G1), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n411), .A2(new_n412), .B1(G77), .B2(new_n248), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n330), .A2(G238), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n221), .B2(new_n333), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n273), .A2(new_n231), .A3(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n292), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n302), .B1(G244), .B2(new_n305), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n421), .B2(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G200), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n321), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n414), .B1(new_n423), .B2(new_n339), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n422), .A2(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n396), .A2(new_n403), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n328), .A2(new_n368), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT75), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n328), .A2(new_n368), .A3(new_n431), .A4(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n330), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n333), .A2(KEYINPUT4), .A3(G244), .A4(new_n329), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n329), .A2(G244), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n284), .B2(new_n285), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n435), .B(new_n436), .C1(new_n438), .C2(KEYINPUT4), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n292), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT5), .B(G41), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n304), .ZN(new_n446));
  INV_X1    g0246(.A(G257), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n442), .A2(new_n304), .A3(G274), .A4(new_n444), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n445), .A2(KEYINPUT76), .A3(G257), .A4(new_n304), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n450), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n292), .B1(new_n444), .B2(new_n442), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT76), .B1(new_n454), .B2(G257), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT77), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n440), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT79), .B1(new_n457), .B2(G179), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n249), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n208), .A2(G33), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n248), .A2(new_n461), .A3(new_n216), .A4(new_n251), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n221), .A2(KEYINPUT6), .A3(G97), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n459), .A2(new_n221), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n467), .B2(KEYINPUT6), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n468), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n275), .B2(new_n221), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n470), .B2(new_n252), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n457), .B2(new_n339), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n473));
  AOI22_X1  g0273(.A1(KEYINPUT77), .A2(new_n473), .B1(new_n439), .B2(new_n292), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT79), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n321), .A4(new_n452), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n458), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n457), .A2(G200), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n440), .A2(G190), .A3(new_n452), .A4(new_n456), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(KEYINPUT78), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(KEYINPUT78), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n471), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n458), .A2(new_n472), .A3(new_n484), .A4(new_n476), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n220), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G238), .B2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n284), .B2(new_n285), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n271), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n292), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n304), .B(G250), .C1(G1), .C2(new_n443), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n304), .A2(G274), .A3(new_n444), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n492), .A2(KEYINPUT81), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n339), .ZN(new_n501));
  AOI21_X1  g0301(.A(G20), .B1(new_n284), .B2(new_n285), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G68), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT19), .B1(new_n342), .B2(G97), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n209), .B1(new_n380), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(KEYINPUT82), .ZN(new_n507));
  NOR3_X1   g0307(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(KEYINPUT82), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n255), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n408), .A2(new_n248), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n408), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(new_n462), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n498), .A2(new_n321), .A3(new_n499), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n501), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n499), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT81), .B1(new_n492), .B2(new_n495), .ZN(new_n520));
  OAI21_X1  g0320(.A(G200), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n498), .A2(G190), .A3(new_n499), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n462), .A2(new_n297), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n514), .A4(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n251), .A2(new_n216), .B1(G20), .B2(new_n490), .ZN(new_n528));
  AOI21_X1  g0328(.A(G20), .B1(G33), .B2(G283), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G33), .B2(new_n459), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n530), .A3(KEYINPUT20), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n490), .A2(G20), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G13), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G1), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g0341(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n490), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT84), .B1(new_n462), .B2(new_n490), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT85), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n533), .A2(new_n534), .B1(new_n539), .B2(new_n537), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n543), .A4(new_n542), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G257), .A2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n222), .B2(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n284), .B2(new_n285), .ZN(new_n553));
  INV_X1    g0353(.A(G303), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n333), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n292), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n445), .A2(G270), .A3(new_n304), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT83), .B1(new_n557), .B2(new_n450), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G169), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n527), .B1(new_n549), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n284), .A2(new_n285), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n551), .ZN(new_n565));
  INV_X1    g0365(.A(new_n555), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n557), .A2(new_n450), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n292), .A2(new_n567), .B1(new_n570), .B2(new_n558), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G190), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n561), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n549), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n545), .A2(new_n548), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(G179), .A3(new_n571), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .A4(new_n561), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n563), .A2(new_n574), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n297), .A2(KEYINPUT22), .A3(G20), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n333), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT86), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n333), .A2(KEYINPUT86), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n502), .A2(G87), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(KEYINPUT22), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT23), .B1(new_n221), .B2(G20), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n221), .A2(KEYINPUT23), .A3(G20), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(new_n589), .B1(new_n491), .B2(new_n209), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT24), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  AOI211_X1 g0393(.A(G20), .B(new_n297), .C1(new_n284), .C2(new_n285), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n593), .B(new_n590), .C1(new_n596), .C2(new_n584), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n252), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT25), .B1(new_n249), .B2(new_n221), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n221), .ZN(new_n602));
  INV_X1    g0402(.A(new_n462), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n601), .A2(new_n602), .B1(G107), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n447), .A2(G1698), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G250), .B2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n284), .B2(new_n285), .ZN(new_n608));
  INV_X1    g0408(.A(G294), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n271), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n292), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n454), .A2(G264), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(new_n450), .A3(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(new_n339), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT87), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(new_n617), .A3(new_n612), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(G179), .A3(new_n450), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n605), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n604), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n598), .B2(new_n252), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n616), .A2(new_n450), .A3(new_n618), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n308), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n613), .A2(new_n354), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n526), .A2(new_n578), .A3(new_n621), .A4(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n434), .A2(new_n486), .A3(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n322), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT18), .B1(new_n630), .B2(new_n291), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n291), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n325), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n425), .A2(new_n426), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n403), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n396), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n311), .B(KEYINPUT17), .Z(new_n638));
  OAI211_X1 g0438(.A(new_n631), .B(new_n633), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n364), .A2(new_n367), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n352), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(G169), .B1(new_n492), .B2(new_n495), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT88), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT88), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n516), .A2(new_n517), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n477), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n496), .A2(G200), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n514), .B2(new_n524), .ZN(new_n650));
  NOR4_X1   g0450(.A1(new_n512), .A2(KEYINPUT89), .A3(new_n513), .A4(new_n523), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n522), .B(new_n648), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n646), .A2(new_n647), .A3(new_n652), .A4(new_n645), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n518), .A2(new_n525), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n478), .B2(new_n485), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n645), .B(new_n653), .C1(new_n655), .C2(new_n647), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n599), .A2(new_n604), .B1(new_n614), .B2(new_n619), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n563), .A2(new_n576), .A3(new_n577), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n626), .B1(new_n308), .B2(new_n624), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n652), .B(new_n645), .C1(new_n605), .C2(new_n661), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n486), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n641), .B1(new_n434), .B2(new_n666), .ZN(G369));
  NAND2_X1  g0467(.A1(new_n539), .A2(new_n209), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n575), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n578), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n563), .A2(new_n576), .A3(new_n577), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n621), .A2(new_n627), .ZN(new_n680));
  INV_X1    g0480(.A(new_n673), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n623), .A2(new_n681), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n680), .A2(new_n682), .B1(new_n621), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n659), .A2(new_n681), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n658), .B2(new_n681), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n212), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n508), .A2(new_n490), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n215), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n697));
  INV_X1    g0497(.A(new_n662), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n658), .B2(new_n659), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n621), .A2(new_n676), .A3(KEYINPUT90), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n697), .A2(new_n698), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n646), .A2(KEYINPUT26), .A3(new_n652), .A4(new_n645), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n655), .B2(KEYINPUT26), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n704), .A3(new_n645), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n696), .B1(new_n705), .B2(new_n681), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n696), .B(new_n681), .C1(new_n656), .C2(new_n663), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n605), .A2(new_n661), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n711), .A2(new_n654), .A3(new_n658), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n697), .A3(new_n578), .A4(new_n681), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n500), .A2(new_n457), .ZN(new_n714));
  INV_X1    g0514(.A(new_n618), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n556), .B(G179), .C1(new_n559), .C2(new_n560), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n617), .B1(new_n611), .B2(new_n612), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n718), .A3(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n474), .A2(new_n498), .A3(new_n452), .A4(new_n499), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n616), .A2(new_n571), .A3(G179), .A4(new_n618), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n571), .A2(G179), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n624), .A2(new_n724), .A3(new_n457), .A4(new_n496), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n719), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n726), .B2(new_n673), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n710), .B1(new_n713), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n709), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n695), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n538), .A2(G20), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G45), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G1), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n690), .A2(KEYINPUT91), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT91), .B1(new_n690), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n679), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n677), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n538), .A2(new_n271), .A3(KEYINPUT93), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT93), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G13), .B2(G33), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n216), .B1(G20), .B2(new_n339), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n564), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n212), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT92), .ZN(new_n755));
  INV_X1    g0555(.A(new_n215), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n443), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n755), .B(new_n757), .C1(new_n443), .C2(new_n241), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n689), .A2(new_n273), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G355), .B1(new_n490), .B2(new_n689), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n752), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n750), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n209), .A2(G179), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n354), .A3(G200), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n763), .A2(new_n765), .B1(new_n766), .B2(new_n554), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n209), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n321), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G329), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n770), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n769), .A2(G20), .A3(G190), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n273), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n209), .B1(new_n772), .B2(G190), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n609), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n767), .A2(new_n775), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n209), .A2(new_n321), .A3(new_n308), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n786));
  INV_X1    g0586(.A(G317), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n783), .A2(new_n354), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n781), .B1(new_n785), .B2(new_n788), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G50), .A2(new_n790), .B1(new_n784), .B2(G68), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n773), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n796), .A2(KEYINPUT32), .B1(new_n297), .B2(new_n766), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n765), .A2(new_n221), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n333), .B1(new_n776), .B2(new_n202), .ZN(new_n800));
  INV_X1    g0600(.A(new_n770), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G77), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n779), .A2(new_n459), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n796), .B2(KEYINPUT32), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n793), .A2(new_n799), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n762), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n761), .A2(new_n806), .A3(new_n740), .ZN(new_n807));
  INV_X1    g0607(.A(new_n749), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n677), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n743), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  AOI22_X1  g0611(.A1(new_n422), .A2(new_n424), .B1(new_n415), .B2(new_n673), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(new_n635), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n635), .A2(new_n681), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n666), .B2(new_n673), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n427), .A2(new_n681), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n656), .B2(new_n663), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n741), .B1(new_n819), .B2(new_n731), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n731), .B2(new_n819), .ZN(new_n821));
  INV_X1    g0621(.A(new_n776), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT96), .B(G143), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n822), .A2(new_n824), .B1(new_n801), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n785), .B2(new_n826), .C1(new_n827), .C2(new_n791), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT34), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(new_n765), .ZN(new_n832));
  INV_X1    g0632(.A(new_n779), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(G68), .B1(new_n833), .B2(G58), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n201), .B2(new_n766), .C1(new_n835), .C2(new_n773), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n830), .A2(new_n831), .A3(new_n753), .A4(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G283), .A2(new_n784), .B1(new_n790), .B2(G303), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n776), .A2(new_n609), .B1(new_n773), .B2(new_n771), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n333), .B(new_n839), .C1(G116), .C2(new_n801), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n765), .A2(new_n297), .ZN(new_n841));
  INV_X1    g0641(.A(new_n766), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n803), .B(new_n841), .C1(G107), .C2(new_n842), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n838), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n750), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n747), .A2(new_n750), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n740), .B1(new_n219), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n815), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n845), .B(new_n847), .C1(new_n848), .C2(new_n748), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n821), .A2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n735), .A2(new_n208), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n396), .A2(new_n403), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n378), .A2(new_n673), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n396), .A2(new_n403), .A3(new_n853), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n815), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n628), .A2(new_n486), .A3(new_n673), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n726), .A2(new_n673), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT31), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n857), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT102), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n857), .B(KEYINPUT102), .C1(new_n858), .C2(new_n863), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(KEYINPUT40), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n671), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n317), .A2(new_n318), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n291), .A2(new_n310), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n323), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT100), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(G68), .A3(new_n288), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(new_n264), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n874), .B(new_n252), .C1(new_n877), .C2(KEYINPUT16), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT16), .B1(new_n876), .B2(new_n264), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT100), .B1(new_n879), .B2(new_n255), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n290), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n671), .B1(new_n881), .B2(new_n314), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n630), .B1(new_n881), .B2(new_n314), .ZN(new_n883));
  INV_X1    g0683(.A(new_n872), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n873), .B1(new_n885), .B2(new_n871), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n327), .A2(KEYINPUT101), .A3(new_n882), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT101), .B1(new_n327), .B2(new_n882), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n886), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n633), .A2(new_n631), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n638), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n873), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n632), .A2(new_n884), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n871), .B1(new_n893), .B2(new_n870), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n891), .A2(new_n870), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT103), .B1(new_n868), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n867), .A2(KEYINPUT40), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n889), .A2(new_n897), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n866), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n896), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n889), .ZN(new_n906));
  INV_X1    g0706(.A(new_n864), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n899), .A2(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n434), .B1(new_n713), .B2(new_n729), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n710), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n818), .A2(new_n814), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n855), .ZN(new_n916));
  INV_X1    g0716(.A(new_n856), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n906), .B1(new_n890), .B2(new_n671), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n902), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n396), .A2(new_n673), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n433), .B1(new_n706), .B2(new_n708), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n641), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n851), .B1(new_n913), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n913), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n468), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n468), .A2(KEYINPUT35), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n216), .A2(new_n209), .A3(new_n490), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT97), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(KEYINPUT97), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n756), .A2(new_n259), .A3(G77), .A4(new_n261), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n201), .A2(G68), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n208), .B(G13), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT98), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT99), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n932), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT104), .ZN(G367));
  OAI21_X1  g0747(.A(new_n751), .B1(new_n212), .B2(new_n515), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n755), .B2(new_n237), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n765), .A2(new_n219), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G68), .B2(new_n833), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n202), .B2(new_n766), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n333), .B1(new_n776), .B2(new_n826), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n770), .A2(new_n201), .B1(new_n773), .B2(new_n827), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n794), .B2(new_n785), .C1(new_n791), .C2(new_n823), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT109), .B1(new_n766), .B2(new_n490), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT46), .Z(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n785), .B2(new_n609), .C1(new_n771), .C2(new_n791), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n776), .A2(new_n554), .B1(new_n773), .B2(new_n787), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G283), .B2(new_n801), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n765), .A2(new_n459), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G107), .B2(new_n833), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n753), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n956), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n740), .B(new_n949), .C1(new_n967), .C2(new_n750), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n650), .A2(new_n651), .A3(new_n681), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n645), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n645), .A3(new_n652), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n749), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n697), .B1(new_n471), .B2(new_n681), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n646), .A2(new_n673), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n686), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT42), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n970), .A2(new_n971), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n621), .B1(new_n974), .B2(new_n975), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n478), .A2(new_n485), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n681), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n979), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT105), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n979), .A2(new_n984), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n980), .B(KEYINPUT43), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n985), .A2(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n986), .B2(new_n985), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n679), .A2(new_n976), .A3(new_n683), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n990), .A2(KEYINPUT106), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT106), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n991), .A2(KEYINPUT106), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n737), .B(KEYINPUT107), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n976), .A2(new_n687), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT45), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n976), .A2(new_n687), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT44), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(new_n684), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n683), .B1(new_n659), .B2(new_n681), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(new_n686), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n678), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n732), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n732), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n690), .B(KEYINPUT41), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n998), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n997), .A2(KEYINPUT108), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT108), .B1(new_n997), .B2(new_n1011), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n973), .B1(new_n1013), .B2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n1008), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1007), .A2(new_n732), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n690), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n759), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n692), .B1(G107), .B2(new_n212), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n692), .B(new_n443), .C1(new_n203), .C2(new_n219), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n246), .B2(G50), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n247), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n234), .B2(G45), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1020), .B1(new_n755), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n741), .B1(new_n1027), .B2(new_n752), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G159), .A2(new_n790), .B1(new_n784), .B2(new_n247), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n515), .A2(new_n779), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n962), .B(new_n1030), .C1(G77), .C2(new_n842), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n770), .A2(new_n203), .B1(new_n773), .B2(new_n826), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G50), .B2(new_n822), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n564), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n766), .A2(new_n609), .B1(new_n779), .B2(new_n763), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT111), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n822), .A2(G317), .B1(new_n801), .B2(G303), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n785), .B2(new_n771), .C1(new_n777), .C2(new_n791), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n1039), .B2(new_n1038), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n765), .A2(new_n490), .B1(new_n773), .B2(new_n789), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n564), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1028), .B1(new_n1047), .B2(new_n750), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n683), .B2(new_n808), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT112), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1018), .B(new_n1050), .C1(new_n1007), .C2(new_n998), .ZN(G393));
  INV_X1    g0851(.A(new_n998), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n974), .A2(new_n749), .A3(new_n975), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n790), .A2(G150), .B1(G159), .B2(new_n822), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT51), .Z(new_n1055));
  NAND2_X1  g0855(.A1(new_n784), .A2(G50), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n770), .A2(new_n246), .B1(new_n773), .B2(new_n823), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n766), .A2(new_n203), .B1(new_n779), .B2(new_n219), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n841), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n564), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n790), .A2(G317), .B1(G311), .B2(new_n822), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n273), .B1(new_n773), .B2(new_n777), .C1(new_n609), .C2(new_n770), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n798), .B1(G116), .B2(new_n833), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n763), .B2(new_n766), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G303), .C2(new_n784), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n762), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n755), .A2(new_n244), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n752), .B1(G97), .B2(new_n689), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n740), .B(new_n1068), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1004), .A2(new_n1052), .B1(new_n1053), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1004), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n690), .B1(new_n1073), .B2(new_n1016), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(G390));
  INV_X1    g0876(.A(new_n918), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n925), .B1(new_n914), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT39), .B1(new_n889), .B2(new_n897), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n902), .A2(new_n924), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n705), .A2(new_n681), .A3(new_n813), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n918), .B1(new_n1084), .B2(new_n814), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n730), .A2(new_n1077), .A3(new_n848), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1082), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1087), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1078), .B1(new_n921), .B2(new_n923), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n747), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n846), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n741), .B1(new_n247), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n785), .A2(new_n221), .B1(new_n459), .B2(new_n770), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n203), .A2(new_n765), .B1(new_n766), .B2(new_n297), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n273), .B1(new_n773), .B2(new_n609), .C1(new_n490), .C2(new_n776), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(G77), .C2(new_n833), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1099), .B(new_n1102), .C1(new_n763), .C2(new_n791), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n790), .A2(G128), .B1(G132), .B2(new_n822), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT116), .ZN(new_n1106));
  INV_X1    g0906(.A(G125), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n333), .B1(new_n773), .B2(new_n1107), .C1(new_n201), .C2(new_n765), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT115), .Z(new_n1109));
  NOR2_X1   g0909(.A1(new_n766), .A2(new_n826), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n770), .A2(new_n1112), .B1(new_n779), .B2(new_n794), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n784), .B2(G137), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1109), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1103), .A2(new_n1104), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1097), .B1(new_n1116), .B2(new_n750), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1094), .A2(new_n1052), .B1(new_n1095), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n433), .A2(new_n730), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n928), .A2(new_n641), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1077), .B1(new_n730), .B2(new_n848), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n914), .B1(new_n1089), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1123), .A2(new_n814), .A3(new_n1084), .A4(new_n1087), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1120), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1088), .A2(new_n1092), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT113), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT113), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1088), .A2(new_n1092), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1125), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n691), .B1(new_n1093), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(KEYINPUT114), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT114), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1118), .B1(new_n1134), .B2(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(KEYINPUT57), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n899), .A2(new_n903), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n710), .B1(new_n908), .B2(new_n909), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n368), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n671), .B1(new_n358), .B2(new_n360), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1139), .A2(new_n1140), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n927), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1150), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n927), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1139), .A2(new_n1140), .A3(new_n1150), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1120), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1138), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1120), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1130), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1138), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n691), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT121), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1163), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1160), .A2(KEYINPUT57), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n690), .C1(new_n1170), .C2(new_n1162), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1155), .A2(new_n747), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n741), .B1(G50), .B2(new_n1096), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n515), .A2(new_n770), .B1(new_n763), .B2(new_n773), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n842), .A2(G77), .B1(new_n833), .B2(G68), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n202), .B2(new_n765), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G107), .C2(new_n822), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n753), .A2(new_n303), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G97), .B2(new_n784), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n490), .C2(new_n791), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT58), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1180), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n766), .A2(new_n1112), .ZN(new_n1188));
  INV_X1    g0988(.A(G128), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n776), .A2(new_n1189), .B1(new_n770), .B2(new_n827), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(G150), .C2(new_n833), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n785), .B2(new_n835), .C1(new_n1107), .C2(new_n791), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT120), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n832), .A2(G159), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n773), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G33), .B(G41), .C1(new_n1198), .C2(G124), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1187), .B1(KEYINPUT58), .B2(new_n1183), .C1(new_n1195), .C2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1175), .B1(new_n1201), .B2(new_n750), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1160), .A2(new_n1052), .B1(new_n1174), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1173), .A2(new_n1203), .ZN(G375));
  INV_X1    g1004(.A(new_n1010), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1124), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1131), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n998), .B1(new_n1124), .B2(new_n1122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n918), .A2(new_n747), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n741), .B1(G68), .B2(new_n1096), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G116), .A2(new_n784), .B1(new_n790), .B2(G294), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n776), .A2(new_n763), .B1(new_n773), .B2(new_n554), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n333), .B(new_n1212), .C1(G107), .C2(new_n801), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n950), .B(new_n1030), .C1(G97), .C2(new_n842), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n766), .A2(new_n794), .B1(new_n779), .B2(new_n201), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n776), .A2(new_n827), .B1(new_n773), .B2(new_n1189), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G150), .C2(new_n801), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n785), .B2(new_n1112), .C1(new_n835), .C2(new_n791), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n564), .B1(new_n202), .B2(new_n765), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT122), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1210), .B1(new_n1222), .B2(new_n750), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1208), .B1(new_n1209), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1207), .A2(new_n1224), .ZN(G381));
  INV_X1    g1025(.A(G387), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1224), .A3(new_n1207), .A4(new_n1227), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1133), .A2(new_n1118), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OR3_X1    g1030(.A1(new_n1228), .A2(G375), .A3(new_n1230), .ZN(G407));
  NAND2_X1  g1031(.A1(new_n672), .A2(G213), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G375), .C2(new_n1234), .ZN(G409));
  OAI211_X1 g1035(.A(G378), .B(new_n1203), .C1(new_n1169), .C2(new_n1172), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n998), .B1(new_n1160), .B2(KEYINPUT123), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(KEYINPUT123), .B2(new_n1160), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1174), .A2(new_n1202), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1161), .A2(new_n1162), .A3(new_n1010), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1229), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1232), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n691), .B1(new_n1245), .B2(new_n1206), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1206), .B2(new_n1245), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1247), .A2(new_n1224), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(G384), .B(KEYINPUT124), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1224), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G2897), .B(new_n1233), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1233), .A2(G2897), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1253), .B(new_n1256), .C1(new_n1248), .C2(new_n1250), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1244), .B2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1243), .A2(new_n1232), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(G387), .B2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G393), .B(new_n810), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(G387), .A2(new_n1266), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1014), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1012), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G390), .B1(new_n1271), .B2(new_n973), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1267), .A2(new_n1268), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1226), .A2(G390), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(new_n1266), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1265), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1233), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1260), .A2(new_n1264), .A3(new_n1278), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1278), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1279), .B2(new_n1258), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1262), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1279), .A2(KEYINPUT62), .A3(new_n1261), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1284), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1282), .B1(new_n1288), .B2(KEYINPUT126), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1287), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT62), .B1(new_n1279), .B2(new_n1261), .ZN(new_n1291));
  OAI211_X1 g1091(.A(KEYINPUT126), .B(new_n1260), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1281), .B1(new_n1289), .B2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1261), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1273), .B(new_n1277), .C1(new_n1254), .C2(new_n1251), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1236), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(G375), .B2(new_n1229), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1297), .B(new_n1299), .ZN(G402));
endmodule


