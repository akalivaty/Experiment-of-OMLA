//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G244), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n215), .A2(G77), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G226), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G68), .B(G77), .ZN(new_n235));
  INV_X1    g0035(.A(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT67), .B(G50), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NOR2_X1   g0043(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n244));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n211), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n250), .A2(new_n252), .B1(G50), .B2(new_n249), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT70), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n212), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(G150), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G50), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n212), .B1(new_n201), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT69), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n247), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT9), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OR3_X1    g0066(.A1(new_n254), .A2(new_n265), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n271), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G226), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G223), .A3(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G222), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n287), .B1(new_n288), .B2(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n270), .A2(KEYINPUT68), .A3(new_n271), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT68), .B1(new_n270), .B2(new_n271), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n281), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G200), .B1(KEYINPUT73), .B2(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(G190), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n244), .B1(new_n268), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  INV_X1    g0102(.A(new_n244), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n266), .A4(new_n267), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n297), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n264), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n255), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n251), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n313), .A2(new_n250), .B1(new_n249), .B2(new_n312), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT16), .ZN(new_n315));
  INV_X1    g0115(.A(G68), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n236), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n317), .B2(new_n201), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n258), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n284), .A2(new_n212), .A3(new_n285), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n285), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT77), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n321), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(KEYINPUT77), .B(new_n316), .C1(new_n324), .C2(new_n325), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n315), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n326), .A2(new_n320), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n247), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n314), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n293), .A2(new_n294), .ZN(new_n335));
  AND2_X1   g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  OAI211_X1 g0137(.A(G226), .B(G1698), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT78), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n286), .A2(new_n340), .A3(G226), .A4(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(G223), .B(new_n289), .C1(new_n336), .C2(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n335), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G232), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n276), .B1(new_n279), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n334), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n349), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n345), .B1(new_n341), .B2(new_n339), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n335), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n333), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT17), .ZN(new_n357));
  OAI21_X1  g0157(.A(G169), .B1(new_n347), .B2(new_n349), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n351), .B(G179), .C1(new_n353), .C2(new_n335), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT18), .B1(new_n333), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n314), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n336), .A2(new_n337), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n212), .ZN(new_n364));
  INV_X1    g0164(.A(new_n325), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n320), .B1(new_n366), .B2(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n326), .A2(new_n327), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT16), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n321), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n246), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n362), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n358), .A2(new_n359), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT79), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n361), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n361), .B2(new_n375), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n357), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(G226), .B(new_n289), .C1(new_n336), .C2(new_n337), .ZN(new_n381));
  OAI211_X1 g0181(.A(G232), .B(G1698), .C1(new_n336), .C2(new_n337), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n295), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n275), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G238), .B1(new_n275), .B2(new_n272), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n385), .B2(new_n388), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT14), .B1(new_n392), .B2(new_n308), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(G169), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT76), .B1(new_n392), .B2(G179), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n390), .A2(new_n391), .A3(new_n397), .A4(new_n306), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n393), .B(new_n395), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n256), .A2(new_n288), .B1(new_n212), .B2(G68), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(KEYINPUT74), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(KEYINPUT74), .B1(G50), .B2(new_n258), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT11), .A3(new_n246), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n249), .A2(G68), .B1(KEYINPUT75), .B2(KEYINPUT12), .ZN(new_n405));
  NAND2_X1  g0205(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(new_n250), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n316), .B1(new_n248), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT11), .B1(new_n403), .B2(new_n246), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n399), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G200), .B1(new_n390), .B2(new_n391), .ZN(new_n417));
  INV_X1    g0217(.A(new_n391), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(G190), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n414), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT15), .B(G87), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n424), .A2(new_n256), .B1(new_n212), .B2(new_n288), .ZN(new_n425));
  INV_X1    g0225(.A(new_n258), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n255), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n247), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT72), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n251), .A2(G77), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n250), .A2(new_n431), .B1(G77), .B2(new_n249), .ZN(new_n432));
  OR3_X1    g0232(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n286), .A2(G238), .A3(G1698), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT71), .B(G107), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n435), .B1(new_n437), .B2(new_n286), .C1(new_n290), .C2(new_n348), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n295), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n387), .A2(new_n215), .B1(new_n275), .B2(new_n272), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(G190), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n433), .A2(new_n434), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n440), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G200), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n433), .A2(new_n434), .B1(new_n308), .B2(new_n443), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n439), .A2(new_n306), .A3(new_n440), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NOR4_X1   g0251(.A1(new_n311), .A2(new_n380), .A3(new_n423), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n286), .A2(new_n212), .A3(G87), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT22), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT22), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n286), .A2(new_n455), .A3(new_n212), .A4(G87), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n458), .A2(G107), .B1(new_n459), .B2(new_n256), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n437), .A2(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(KEYINPUT23), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n457), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n457), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n246), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n247), .B(new_n249), .C1(G1), .C2(new_n283), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n249), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT25), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(KEYINPUT25), .A3(new_n470), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n468), .A2(G107), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n286), .A2(G257), .A3(G1698), .ZN(new_n475));
  OAI211_X1 g0275(.A(G250), .B(new_n289), .C1(new_n336), .C2(new_n337), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n274), .A2(G1), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT5), .B(G41), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n386), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n478), .A2(new_n295), .B1(G264), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n272), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(G190), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G200), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n466), .A2(new_n474), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n308), .B1(new_n482), .B2(new_n484), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(G179), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n466), .A2(new_n474), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n488), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n469), .A2(new_n459), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n467), .B2(new_n459), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n245), .A2(new_n211), .B1(G20), .B2(new_n459), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n212), .C1(G33), .C2(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n499), .A2(KEYINPUT20), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT20), .B1(new_n499), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(KEYINPUT21), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n481), .A2(G270), .B1(new_n483), .B2(new_n272), .ZN(new_n511));
  OAI211_X1 g0311(.A(G264), .B(G1698), .C1(new_n336), .C2(new_n337), .ZN(new_n512));
  OAI211_X1 g0312(.A(G257), .B(new_n289), .C1(new_n336), .C2(new_n337), .ZN(new_n513));
  XOR2_X1   g0313(.A(KEYINPUT81), .B(G303), .Z(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n286), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n295), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n507), .A2(G169), .A3(new_n510), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n517), .ZN(new_n519));
  OAI21_X1  g0319(.A(G169), .B1(new_n498), .B2(new_n505), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n509), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n511), .A2(G179), .A3(new_n516), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n522), .A2(new_n506), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n518), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(G190), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n517), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n506), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT83), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n525), .A2(new_n529), .A3(new_n506), .A4(new_n526), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n524), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n501), .A2(new_n470), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n470), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT80), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT6), .A2(G97), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n436), .B1(new_n364), .B2(new_n365), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n247), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n249), .A2(G97), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n468), .B2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  INV_X1    g0348(.A(G244), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n286), .A2(new_n289), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n284), .B2(new_n285), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n500), .C1(KEYINPUT4), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n286), .A2(G250), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n289), .B1(new_n554), .B2(KEYINPUT4), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n295), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n481), .A2(G257), .B1(new_n483), .B2(new_n272), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n547), .B(new_n559), .C1(new_n352), .C2(new_n558), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n541), .A2(new_n542), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n545), .B1(new_n561), .B2(new_n247), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n558), .A2(new_n308), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n306), .A3(new_n557), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n286), .A2(G238), .A3(new_n289), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(G1698), .C1(new_n336), .C2(new_n337), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G116), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n295), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n248), .A2(new_n269), .A3(G45), .ZN(new_n572));
  INV_X1    g0372(.A(G250), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n274), .B2(G1), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n277), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G169), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n575), .ZN(new_n577));
  AOI211_X1 g0377(.A(G179), .B(new_n577), .C1(new_n570), .C2(new_n295), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n424), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n249), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n212), .B1(new_n383), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n501), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n436), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n286), .A2(new_n212), .A3(G68), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n582), .B1(new_n256), .B2(new_n501), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n581), .B1(new_n589), .B2(new_n246), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n424), .B2(new_n467), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n579), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n577), .B1(new_n570), .B2(new_n295), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n593), .A2(new_n334), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n468), .A2(G87), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n590), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n566), .A2(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n452), .A2(new_n496), .A3(new_n531), .A4(new_n599), .ZN(G372));
  NOR2_X1   g0400(.A1(new_n593), .A2(new_n334), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n590), .A2(new_n596), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n595), .B1(new_n579), .B2(new_n591), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n466), .A2(new_n474), .A3(new_n485), .A4(new_n487), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n560), .A3(new_n605), .A4(new_n565), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n493), .A2(new_n492), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n495), .B1(new_n608), .B2(new_n490), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n521), .A2(new_n523), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n518), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n607), .A2(new_n611), .B1(new_n591), .B2(new_n579), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n564), .B1(new_n543), .B2(new_n546), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n481), .A2(G257), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n484), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n363), .A2(new_n573), .ZN(new_n617));
  OAI21_X1  g0417(.A(G1698), .B1(new_n617), .B2(new_n548), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n286), .A2(G244), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(new_n548), .B1(G33), .B2(G283), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n620), .A3(new_n551), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n616), .B1(new_n621), .B2(new_n295), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G169), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n613), .B1(new_n614), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT85), .A4(new_n564), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n604), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT86), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n614), .A2(new_n623), .ZN(new_n629));
  XNOR2_X1  g0429(.A(KEYINPUT87), .B(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n604), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT88), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT88), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n604), .A2(new_n629), .A3(new_n634), .A4(new_n631), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT86), .B1(new_n626), .B2(new_n627), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n612), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n452), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT89), .Z(new_n640));
  INV_X1    g0440(.A(new_n310), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n333), .A2(new_n360), .A3(KEYINPUT18), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n374), .B1(new_n372), .B2(new_n373), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n357), .A2(new_n422), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n449), .B1(new_n415), .B2(new_n399), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n641), .B1(new_n647), .B2(new_n305), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n640), .A2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n248), .A2(new_n212), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n506), .A2(new_n656), .ZN(new_n657));
  MUX2_X1   g0457(.A(new_n531), .B(new_n524), .S(new_n657), .Z(new_n658));
  XNOR2_X1  g0458(.A(KEYINPUT90), .B(G330), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n495), .A2(new_n655), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n496), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n609), .B2(new_n656), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n494), .A2(new_n495), .A3(new_n656), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n524), .A2(new_n656), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n496), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n206), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n436), .A2(G116), .A3(new_n585), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n209), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n630), .B1(new_n598), .B2(new_n565), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n624), .A2(new_n604), .A3(new_n625), .A4(KEYINPUT26), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n680), .B(new_n630), .C1(new_n598), .C2(new_n565), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n607), .A2(KEYINPUT93), .A3(new_n611), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT93), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n524), .B1(new_n494), .B2(new_n495), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n606), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n682), .A2(new_n683), .A3(new_n686), .A4(new_n592), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .A3(new_n656), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n626), .A2(new_n627), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT86), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n628), .A3(new_n633), .A4(new_n635), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n655), .B1(new_n692), .B2(new_n612), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n688), .B1(new_n693), .B2(KEYINPUT29), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n496), .A2(new_n599), .A3(new_n531), .A4(new_n656), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n482), .A2(new_n593), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n558), .A2(new_n696), .A3(new_n522), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT91), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT30), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n696), .A2(new_n522), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT91), .B(new_n700), .C1(new_n701), .C2(new_n558), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n519), .A2(G179), .A3(new_n593), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n486), .A3(new_n558), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n699), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n655), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n695), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n660), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n694), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n676), .B1(new_n713), .B2(G1), .ZN(G364));
  AND2_X1   g0514(.A1(new_n212), .A2(G13), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n248), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n671), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n661), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n660), .B2(new_n658), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n286), .A2(new_n206), .ZN(new_n721));
  INV_X1    g0521(.A(G355), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n721), .A2(new_n722), .B1(G116), .B2(new_n206), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n363), .A2(new_n206), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n274), .B2(new_n210), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n239), .A2(G45), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n211), .B1(G20), .B2(new_n308), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n718), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n212), .A2(new_n306), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G200), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT95), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT33), .B(G317), .ZN(new_n741));
  INV_X1    g0541(.A(new_n737), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n352), .A3(G200), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(new_n741), .B1(G322), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n286), .B1(new_n746), .B2(G311), .ZN(new_n747));
  INV_X1    g0547(.A(G283), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n212), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n352), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n747), .B1(new_n748), .B2(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  OR3_X1    g0553(.A1(KEYINPUT96), .A2(G179), .A3(G200), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT96), .B1(G179), .B2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n212), .A2(G190), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n753), .B1(G329), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n739), .A2(new_n352), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n352), .B1(new_n754), .B2(new_n755), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n212), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n760), .A2(G326), .B1(G294), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n745), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n584), .A2(new_n752), .B1(new_n750), .B2(new_n470), .ZN(new_n766));
  INV_X1    g0566(.A(new_n746), .ZN(new_n767));
  INV_X1    g0567(.A(new_n743), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n286), .B1(new_n767), .B2(new_n288), .C1(new_n236), .C2(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n766), .B(new_n769), .C1(new_n740), .C2(G68), .ZN(new_n770));
  INV_X1    g0570(.A(new_n758), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(KEYINPUT32), .B1(G97), .B2(new_n763), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT32), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(new_n773), .B1(new_n760), .B2(G50), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n770), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n765), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n736), .B1(new_n779), .B2(new_n733), .ZN(new_n780));
  INV_X1    g0580(.A(new_n732), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n658), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n720), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  NAND2_X1  g0584(.A1(new_n433), .A2(new_n434), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n442), .A2(new_n444), .B1(new_n785), .B2(new_n655), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n449), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n447), .A2(new_n448), .A3(new_n656), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n693), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT100), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n450), .A2(new_n656), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n638), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n718), .B1(new_n795), .B2(new_n711), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n711), .B2(new_n795), .ZN(new_n797));
  INV_X1    g0597(.A(new_n718), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n733), .A2(new_n730), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n288), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G143), .A2(new_n743), .B1(new_n746), .B2(G159), .ZN(new_n801));
  INV_X1    g0601(.A(new_n760), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G150), .B2(new_n740), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT34), .Z(new_n806));
  NOR2_X1   g0606(.A1(new_n762), .A2(new_n236), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n363), .B1(new_n758), .B2(G132), .ZN(new_n808));
  INV_X1    g0608(.A(new_n750), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G68), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n260), .B2(new_n752), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n811), .B2(KEYINPUT99), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n807), .B(new_n812), .C1(KEYINPUT99), .C2(new_n811), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n740), .B(KEYINPUT98), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G283), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n802), .A2(new_n751), .B1(new_n762), .B2(new_n501), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n771), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n363), .B1(new_n767), .B2(new_n459), .C1(new_n820), .C2(new_n768), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n584), .A2(new_n750), .B1(new_n752), .B2(new_n470), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n817), .A2(new_n819), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n806), .A2(new_n813), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n733), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n800), .B1(new_n731), .B2(new_n789), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n797), .A2(new_n826), .ZN(G384));
  OR2_X1    g0627(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n828), .A2(G116), .A3(new_n213), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT36), .Z(new_n831));
  OR3_X1    g0631(.A1(new_n209), .A2(new_n288), .A3(new_n317), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n260), .A2(G68), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n248), .B(G13), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n653), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n644), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n415), .B(new_n655), .C1(new_n399), .C2(new_n421), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n414), .A2(new_n656), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n421), .B(new_n840), .C1(new_n399), .C2(new_n415), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n788), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n794), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n315), .B1(new_n326), .B2(new_n320), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(KEYINPUT101), .A3(new_n246), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n370), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT101), .B1(new_n846), .B2(new_n246), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n362), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n836), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT79), .B1(new_n642), .B2(new_n643), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n377), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n853), .B2(new_n357), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n850), .A2(new_n373), .B1(new_n333), .B2(new_n355), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n851), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n330), .A2(new_n332), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n858), .A2(new_n355), .A3(new_n362), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n858), .A2(new_n362), .B1(new_n358), .B2(new_n359), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n372), .A2(new_n836), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n855), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n372), .A2(new_n373), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n865), .A2(new_n863), .A3(new_n855), .A4(new_n356), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n857), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n845), .B1(new_n854), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n851), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n380), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n857), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n837), .B1(new_n844), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n854), .A2(new_n868), .A3(new_n845), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n861), .A2(new_n863), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n873), .B2(new_n874), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n357), .A2(new_n644), .ZN(new_n884));
  INV_X1    g0684(.A(new_n863), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n879), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n416), .A2(new_n655), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n869), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n878), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n452), .B(new_n688), .C1(new_n693), .C2(KEYINPUT29), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n648), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n892), .B(new_n894), .Z(new_n895));
  OAI21_X1  g0695(.A(new_n789), .B1(new_n839), .B2(new_n841), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n695), .A2(new_n709), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n706), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n705), .A2(KEYINPUT103), .A3(new_n655), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n707), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n896), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n880), .B2(new_n887), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n843), .B1(new_n786), .B2(new_n449), .ZN(new_n905));
  INV_X1    g0705(.A(new_n840), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n416), .A2(new_n422), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n838), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n705), .A2(KEYINPUT103), .A3(new_n655), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT103), .B1(new_n705), .B2(new_n655), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT31), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n695), .A2(new_n709), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n904), .B(new_n908), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n903), .A2(KEYINPUT40), .B1(new_n914), .B2(new_n877), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n897), .A2(new_n901), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n452), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n895), .B1(new_n659), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n248), .B2(new_n715), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n895), .A2(new_n659), .A3(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n835), .B1(new_n920), .B2(new_n921), .ZN(G367));
  NAND2_X1  g0722(.A1(new_n602), .A2(new_n655), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n604), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n592), .B2(new_n923), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(new_n781), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n725), .A2(new_n233), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n735), .B1(new_n670), .B2(new_n580), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n798), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n815), .A2(G159), .B1(G50), .B2(new_n746), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n762), .A2(new_n316), .ZN(new_n933));
  INV_X1    g0733(.A(G150), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n286), .B1(new_n236), .B2(new_n752), .C1(new_n768), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G77), .B2(new_n809), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n803), .B2(new_n771), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n933), .B(new_n937), .C1(G143), .C2(new_n760), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n932), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT108), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n752), .A2(new_n459), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n814), .C2(new_n820), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n802), .A2(new_n818), .B1(new_n762), .B2(new_n437), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n363), .B1(new_n767), .B2(new_n748), .C1(new_n514), .C2(new_n768), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n501), .B2(new_n750), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n948), .B(new_n951), .C1(G317), .C2(new_n758), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n940), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT47), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n825), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n955), .A2(new_n956), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n926), .B(new_n929), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n668), .A2(new_n666), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n560), .B(new_n565), .C1(new_n547), .C2(new_n656), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n629), .A2(new_n655), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n961), .A2(new_n965), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT105), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT44), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(new_n661), .A3(new_n664), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n967), .B(new_n665), .C1(new_n972), .C2(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n668), .B1(new_n664), .B2(new_n667), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n661), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n713), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n713), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n671), .B(KEYINPUT41), .Z(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n717), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n964), .A2(new_n496), .A3(new_n667), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n565), .B1(new_n962), .B2(new_n609), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n656), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT104), .Z(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n665), .A2(new_n965), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n960), .B1(new_n984), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT109), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT109), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(G387));
  OR2_X1    g0802(.A1(new_n664), .A2(new_n781), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n673), .A2(new_n721), .B1(G107), .B2(new_n206), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT110), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n230), .A2(G45), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n673), .ZN(new_n1007));
  AOI211_X1 g0807(.A(G45), .B(new_n1007), .C1(G68), .C2(G77), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n255), .A2(G50), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n726), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1005), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n718), .B1(new_n1012), .B2(new_n735), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n286), .B1(new_n767), .B2(new_n316), .C1(new_n260), .C2(new_n768), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G97), .B2(new_n809), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n752), .A2(new_n288), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT111), .B(G150), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(new_n758), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT112), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n762), .A2(new_n424), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G159), .A2(new_n760), .B1(new_n740), .B2(new_n312), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1015), .A2(new_n1019), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n760), .A2(G322), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n743), .A2(G317), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n514), .C2(new_n767), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n814), .B2(new_n818), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n762), .A2(new_n748), .B1(new_n820), .B2(new_n752), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(KEYINPUT49), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n758), .A2(G326), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n286), .B1(new_n809), .B2(G116), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT49), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1023), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1013), .B1(new_n1038), .B2(new_n733), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n979), .A2(new_n717), .B1(new_n1003), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n980), .A2(new_n671), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n713), .A2(new_n979), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  NAND3_X1  g0843(.A1(new_n975), .A2(new_n717), .A3(new_n976), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n734), .B1(new_n501), .B2(new_n206), .C1(new_n726), .C2(new_n242), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n718), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n762), .A2(new_n288), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n363), .B1(new_n746), .B2(new_n312), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n316), .B2(new_n752), .C1(new_n584), .C2(new_n750), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(G143), .C2(new_n758), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n760), .A2(G150), .B1(G159), .B2(new_n743), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1052));
  XNOR2_X1  g0852(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1053), .C1(new_n260), .C2(new_n814), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n760), .A2(G317), .B1(G311), .B2(new_n743), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  NOR2_X1   g0857(.A1(new_n762), .A2(new_n459), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n286), .B1(new_n746), .B2(G294), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n470), .B2(new_n750), .C1(new_n748), .C2(new_n752), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(G322), .C2(new_n758), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1057), .B(new_n1061), .C1(new_n514), .C2(new_n814), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1055), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1046), .B1(new_n1064), .B2(new_n733), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n781), .B2(new_n964), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1044), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT115), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n977), .A2(new_n980), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n977), .A2(new_n980), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n671), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(G390));
  NAND2_X1  g0872(.A1(new_n888), .A2(new_n890), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n842), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n792), .B1(new_n692), .B2(new_n612), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n788), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n889), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n787), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n687), .A2(new_n656), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n843), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1074), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n864), .A2(new_n867), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n863), .B1(new_n357), .B2(new_n644), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n845), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n889), .B1(new_n876), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1073), .A2(new_n1078), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n916), .A2(G330), .A3(new_n908), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT116), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT116), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1088), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n888), .A2(new_n890), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1077), .B1(new_n880), .B2(new_n887), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1090), .B(new_n1091), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1074), .A2(new_n660), .A3(new_n710), .A4(new_n789), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1089), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n452), .A2(G330), .A3(new_n916), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n893), .A2(new_n648), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n916), .A2(G330), .A3(new_n789), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n842), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1102), .A2(new_n843), .A3(new_n1080), .A4(new_n1096), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n842), .B1(new_n711), .B2(new_n905), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1088), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1075), .B2(new_n788), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1100), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1089), .A2(new_n1095), .A3(new_n1097), .A4(new_n1107), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n671), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n798), .B1(new_n255), .B2(new_n799), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n810), .B1(new_n768), .B2(new_n459), .C1(new_n501), .C2(new_n767), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1047), .B(new_n1113), .C1(G294), .C2(new_n758), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n752), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n286), .B1(new_n1115), .B2(G87), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n802), .A2(new_n748), .B1(new_n1116), .B2(KEYINPUT117), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(KEYINPUT117), .B2(new_n1116), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1114), .B(new_n1118), .C1(new_n437), .C2(new_n814), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n814), .A2(new_n803), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n363), .B1(new_n743), .B2(G132), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1121), .B1(new_n260), .B2(new_n750), .C1(new_n767), .C2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G125), .B2(new_n758), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n760), .A2(G128), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1115), .A2(new_n1017), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G159), .B2(new_n763), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1124), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1119), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n733), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1112), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1073), .B2(new_n730), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1089), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n717), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1111), .A2(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(G330), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n914), .A2(new_n877), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n892), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n891), .B(new_n878), .C1(new_n915), .C2(new_n1140), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n264), .A2(new_n836), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT120), .Z(new_n1147));
  OR2_X1    g0947(.A1(new_n311), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n311), .A2(new_n1147), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1149), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1144), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n717), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n286), .A2(G41), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(G33), .A2(G41), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1157), .A2(G50), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n933), .B1(new_n740), .B2(G97), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n459), .B2(new_n802), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n767), .B2(new_n424), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G107), .B2(new_n743), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n236), .B2(new_n750), .C1(new_n288), .C2(new_n752), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1161), .B(new_n1164), .C1(G283), .C2(new_n758), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1159), .B1(new_n1165), .B2(KEYINPUT58), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT119), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G128), .A2(new_n743), .B1(new_n746), .B2(G137), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n752), .B2(new_n1122), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n740), .B2(G132), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n760), .A2(G125), .B1(G150), .B2(new_n763), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n758), .A2(G124), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n1158), .C1(new_n772), .C2(new_n750), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1172), .B2(KEYINPUT59), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1165), .A2(KEYINPUT58), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n825), .B1(new_n1167), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n798), .B(new_n1178), .C1(new_n260), .C2(new_n799), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1153), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n731), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1100), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1110), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n671), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1110), .A2(new_n1184), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1180), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1144), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1187), .B2(new_n1193), .ZN(G375));
  NAND2_X1  g0994(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n717), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n842), .A2(new_n730), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n733), .A2(G68), .A3(new_n730), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n288), .A2(new_n750), .B1(new_n752), .B2(new_n501), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n363), .B1(new_n768), .B2(new_n748), .C1(new_n437), .C2(new_n767), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G303), .C2(new_n758), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1020), .B1(new_n760), .B2(G294), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n459), .C2(new_n814), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT122), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n236), .A2(new_n750), .B1(new_n752), .B2(new_n772), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n286), .B1(new_n767), .B2(new_n934), .C1(new_n803), .C2(new_n768), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G128), .C2(new_n758), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n760), .A2(G132), .B1(G50), .B2(new_n763), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n814), .C2(new_n1122), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n798), .B(new_n1198), .C1(new_n1212), .C2(new_n733), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1196), .A2(KEYINPUT121), .B1(new_n1197), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT121), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1195), .A2(new_n1215), .A3(new_n717), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1100), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1108), .A2(new_n983), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(G381));
  OR2_X1    g1022(.A1(G393), .A2(G396), .ZN(new_n1223));
  OR4_X1    g1023(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1223), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G387), .A2(new_n1224), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1025(.A1(new_n654), .A2(G213), .ZN(new_n1226));
  OR3_X1    g1026(.A1(G375), .A2(G378), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G407), .A2(new_n1227), .A3(G213), .ZN(G409));
  INV_X1    g1028(.A(new_n998), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1229), .A2(G390), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(G390), .B(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1231), .B1(new_n1233), .B2(new_n1001), .ZN(new_n1234));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(new_n998), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1229), .A2(G390), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1223), .B(new_n1230), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1183), .C1(new_n1187), .C2(new_n1193), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1188), .A2(new_n1192), .A3(new_n983), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1111), .B(new_n1138), .C1(new_n1243), .C2(new_n1182), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(new_n1226), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1220), .A2(KEYINPUT60), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1220), .A2(KEYINPUT60), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n671), .B(new_n1108), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1219), .A2(G384), .A3(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT123), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1241), .B1(new_n1246), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1245), .A2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1242), .A2(new_n1244), .A3(KEYINPUT124), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n1226), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1257), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1261), .A2(new_n1226), .A3(new_n1263), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n654), .A2(G213), .A3(G2897), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1256), .B(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1259), .B(new_n1265), .C1(new_n1266), .C2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1240), .B1(new_n1268), .B2(new_n1246), .ZN(new_n1270));
  AND4_X1   g1070(.A1(KEYINPUT62), .A2(new_n1262), .A3(new_n1226), .A4(new_n1245), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1264), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1272), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1270), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1269), .B1(new_n1277), .B2(new_n1239), .ZN(G405));
  NAND2_X1  g1078(.A1(new_n1239), .A2(new_n1256), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1234), .A2(new_n1262), .A3(new_n1238), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT127), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G375), .B(G378), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1279), .A2(new_n1284), .A3(new_n1280), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1283), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(G402));
endmodule


