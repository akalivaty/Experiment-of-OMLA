

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U556 ( .A1(n727), .A2(n971), .ZN(n685) );
  AND2_X1 U557 ( .A1(G160), .A2(G40), .ZN(n771) );
  NOR2_X1 U558 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X2 U559 ( .A1(n532), .A2(n531), .ZN(n883) );
  OR2_X1 U560 ( .A1(n894), .A2(n694), .ZN(n695) );
  NOR2_X1 U561 ( .A1(G1966), .A2(n763), .ZN(n741) );
  NOR2_X1 U562 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U563 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U564 ( .A(n770), .B(KEYINPUT99), .ZN(n803) );
  AND2_X1 U565 ( .A1(n541), .A2(n540), .ZN(G160) );
  NOR2_X2 U566 ( .A1(n531), .A2(n532), .ZN(n570) );
  NOR2_X1 U567 ( .A1(n763), .A2(n760), .ZN(n521) );
  NAND2_X4 U568 ( .A1(n773), .A2(n771), .ZN(n727) );
  NOR2_X1 U569 ( .A1(n802), .A2(n523), .ZN(n522) );
  AND2_X1 U570 ( .A1(n1006), .A2(n814), .ZN(n523) );
  AND2_X1 U571 ( .A1(n572), .A2(G137), .ZN(n524) );
  AND2_X1 U572 ( .A1(n534), .A2(n533), .ZN(n525) );
  AND2_X1 U573 ( .A1(n727), .A2(G1341), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n727), .B(KEYINPUT87), .ZN(n697) );
  AND2_X1 U575 ( .A1(n687), .A2(n686), .ZN(n694) );
  XNOR2_X1 U576 ( .A(n737), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U577 ( .A1(G8), .A2(n727), .ZN(n763) );
  XNOR2_X1 U578 ( .A(KEYINPUT13), .B(KEYINPUT67), .ZN(n587) );
  NOR2_X1 U579 ( .A1(n632), .A2(n547), .ZN(n643) );
  NOR2_X1 U580 ( .A1(n632), .A2(G651), .ZN(n647) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n548), .Z(n646) );
  NOR2_X1 U582 ( .A1(n539), .A2(n524), .ZN(n540) );
  XNOR2_X2 U583 ( .A(G2104), .B(KEYINPUT64), .ZN(n531) );
  INV_X1 U584 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G126), .A2(n570), .ZN(n528) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n878) );
  NAND2_X1 U587 ( .A1(G114), .A2(n878), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U589 ( .A(n529), .B(KEYINPUT83), .ZN(n535) );
  NOR2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT17), .B(n530), .Z(n572) );
  NAND2_X1 U592 ( .A1(n572), .A2(G138), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n883), .A2(G102), .ZN(n533) );
  AND2_X2 U594 ( .A1(n535), .A2(n525), .ZN(G164) );
  NAND2_X1 U595 ( .A1(G101), .A2(n883), .ZN(n536) );
  XOR2_X1 U596 ( .A(n536), .B(KEYINPUT23), .Z(n541) );
  NAND2_X1 U597 ( .A1(G125), .A2(n570), .ZN(n538) );
  NAND2_X1 U598 ( .A1(G113), .A2(n878), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT0), .B(G543), .Z(n632) );
  INV_X1 U601 ( .A(G651), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n643), .A2(G76), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT70), .B(n542), .ZN(n545) );
  NOR2_X1 U604 ( .A1(G543), .A2(G651), .ZN(n650) );
  NAND2_X1 U605 ( .A1(n650), .A2(G89), .ZN(n543) );
  XNOR2_X1 U606 ( .A(KEYINPUT4), .B(n543), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n546), .B(KEYINPUT5), .ZN(n554) );
  NOR2_X1 U609 ( .A1(G543), .A2(n547), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n646), .A2(G63), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT71), .B(n549), .Z(n551) );
  NAND2_X1 U612 ( .A1(n647), .A2(G51), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G60), .A2(n646), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G47), .A2(n647), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G85), .A2(n650), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G72), .A2(n643), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  OR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(G290) );
  NAND2_X1 U625 ( .A1(G64), .A2(n646), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G52), .A2(n647), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n643), .A2(G77), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT65), .B(n564), .Z(n566) );
  NAND2_X1 U630 ( .A1(n650), .A2(G90), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(G171) );
  AND2_X1 U634 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U635 ( .A1(G123), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT18), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G99), .A2(n883), .ZN(n574) );
  BUF_X1 U638 ( .A(n572), .Z(n881) );
  NAND2_X1 U639 ( .A1(G135), .A2(n881), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G111), .A2(n878), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT73), .B(n575), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n931) );
  XNOR2_X1 U645 ( .A(G2096), .B(n931), .ZN(n580) );
  OR2_X1 U646 ( .A1(G2100), .A2(n580), .ZN(G156) );
  INV_X1 U647 ( .A(G860), .ZN(n613) );
  NAND2_X1 U648 ( .A1(n646), .A2(G56), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n581), .B(KEYINPUT14), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G43), .A2(n647), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n650), .A2(G81), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G68), .A2(n643), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT68), .B(n591), .Z(n684) );
  BUF_X1 U657 ( .A(n684), .Z(n998) );
  OR2_X1 U658 ( .A1(n613), .A2(n998), .ZN(G153) );
  INV_X1 U659 ( .A(G132), .ZN(G219) );
  INV_X1 U660 ( .A(G82), .ZN(G220) );
  INV_X1 U661 ( .A(G120), .ZN(G236) );
  INV_X1 U662 ( .A(G69), .ZN(G235) );
  INV_X1 U663 ( .A(G108), .ZN(G238) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U666 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n594) );
  INV_X1 U667 ( .A(G223), .ZN(n820) );
  NAND2_X1 U668 ( .A1(G567), .A2(n820), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n594), .B(n593), .ZN(G234) );
  INV_X1 U670 ( .A(G868), .ZN(n664) );
  NOR2_X1 U671 ( .A1(n664), .A2(G171), .ZN(n595) );
  XNOR2_X1 U672 ( .A(n595), .B(KEYINPUT69), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G66), .A2(n646), .ZN(n597) );
  NAND2_X1 U674 ( .A1(G54), .A2(n647), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G92), .A2(n650), .ZN(n599) );
  NAND2_X1 U677 ( .A1(G79), .A2(n643), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT15), .B(n602), .Z(n894) );
  INV_X1 U681 ( .A(n894), .ZN(n1007) );
  NAND2_X1 U682 ( .A1(n664), .A2(n1007), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U684 ( .A1(G65), .A2(n646), .ZN(n606) );
  NAND2_X1 U685 ( .A1(G53), .A2(n647), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G91), .A2(n650), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G78), .A2(n643), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n1001) );
  INV_X1 U691 ( .A(n1001), .ZN(G299) );
  NOR2_X1 U692 ( .A1(G286), .A2(n664), .ZN(n612) );
  NOR2_X1 U693 ( .A1(G868), .A2(G299), .ZN(n611) );
  NOR2_X1 U694 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U695 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n614), .A2(n894), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(KEYINPUT16), .ZN(n616) );
  XNOR2_X1 U698 ( .A(KEYINPUT72), .B(n616), .ZN(G148) );
  NOR2_X1 U699 ( .A1(n998), .A2(G868), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G868), .A2(n894), .ZN(n617) );
  NOR2_X1 U701 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U703 ( .A1(G559), .A2(n894), .ZN(n620) );
  XNOR2_X1 U704 ( .A(n620), .B(n998), .ZN(n662) );
  NOR2_X1 U705 ( .A1(G860), .A2(n662), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G93), .A2(n650), .ZN(n622) );
  NAND2_X1 U707 ( .A1(G80), .A2(n643), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U709 ( .A(KEYINPUT74), .B(n623), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G67), .A2(n646), .ZN(n625) );
  NAND2_X1 U711 ( .A1(G55), .A2(n647), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n665) );
  XOR2_X1 U714 ( .A(n628), .B(n665), .Z(G145) );
  NAND2_X1 U715 ( .A1(G49), .A2(n647), .ZN(n630) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U717 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n646), .A2(n631), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G75), .A2(n643), .ZN(n635) );
  XNOR2_X1 U722 ( .A(n635), .B(KEYINPUT78), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G50), .A2(n647), .ZN(n637) );
  NAND2_X1 U724 ( .A1(G88), .A2(n650), .ZN(n636) );
  NAND2_X1 U725 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U726 ( .A1(G62), .A2(n646), .ZN(n638) );
  XNOR2_X1 U727 ( .A(KEYINPUT77), .B(n638), .ZN(n639) );
  NOR2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(G303) );
  INV_X1 U730 ( .A(G303), .ZN(G166) );
  NAND2_X1 U731 ( .A1(n643), .A2(G73), .ZN(n645) );
  XNOR2_X1 U732 ( .A(KEYINPUT76), .B(KEYINPUT2), .ZN(n644) );
  XNOR2_X1 U733 ( .A(n645), .B(n644), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G61), .A2(n646), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G48), .A2(n647), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G86), .A2(n650), .ZN(n651) );
  XNOR2_X1 U738 ( .A(KEYINPUT75), .B(n651), .ZN(n652) );
  NOR2_X1 U739 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(G305) );
  XNOR2_X1 U741 ( .A(n1001), .B(G288), .ZN(n661) );
  XNOR2_X1 U742 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n657) );
  XOR2_X1 U743 ( .A(G290), .B(n665), .Z(n656) );
  XNOR2_X1 U744 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U745 ( .A(G166), .B(n658), .ZN(n659) );
  XNOR2_X1 U746 ( .A(n659), .B(G305), .ZN(n660) );
  XNOR2_X1 U747 ( .A(n661), .B(n660), .ZN(n893) );
  XOR2_X1 U748 ( .A(n893), .B(n662), .Z(n663) );
  NOR2_X1 U749 ( .A1(n664), .A2(n663), .ZN(n667) );
  NOR2_X1 U750 ( .A1(G868), .A2(n665), .ZN(n666) );
  NOR2_X1 U751 ( .A1(n667), .A2(n666), .ZN(G295) );
  XOR2_X1 U752 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n669) );
  NAND2_X1 U753 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G235), .A2(G236), .ZN(n673) );
  XNOR2_X1 U760 ( .A(n673), .B(KEYINPUT81), .ZN(n674) );
  NOR2_X1 U761 ( .A1(G238), .A2(n674), .ZN(n675) );
  NAND2_X1 U762 ( .A1(G57), .A2(n675), .ZN(n824) );
  NAND2_X1 U763 ( .A1(G567), .A2(n824), .ZN(n680) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U766 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U767 ( .A1(G96), .A2(n678), .ZN(n825) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n825), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U770 ( .A(KEYINPUT82), .B(n681), .Z(G319) );
  INV_X1 U771 ( .A(G319), .ZN(n683) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n682) );
  NOR2_X1 U773 ( .A1(n683), .A2(n682), .ZN(n823) );
  NAND2_X1 U774 ( .A1(n823), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G171), .ZN(G301) );
  NOR2_X2 U776 ( .A1(G164), .A2(G1384), .ZN(n773) );
  NOR2_X1 U777 ( .A1(n684), .A2(n526), .ZN(n687) );
  INV_X1 U778 ( .A(G1996), .ZN(n971) );
  XOR2_X1 U779 ( .A(n685), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U780 ( .A1(n894), .A2(n694), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n697), .A2(G2067), .ZN(n688) );
  XNOR2_X1 U782 ( .A(n688), .B(KEYINPUT90), .ZN(n690) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n727), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U785 ( .A(KEYINPUT91), .B(n691), .Z(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n703) );
  XOR2_X1 U788 ( .A(KEYINPUT27), .B(KEYINPUT89), .Z(n699) );
  NAND2_X1 U789 ( .A1(G2072), .A2(n697), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n699), .B(n698), .ZN(n701) );
  XOR2_X1 U791 ( .A(KEYINPUT87), .B(n727), .Z(n710) );
  AND2_X1 U792 ( .A1(n710), .A2(G1956), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n704), .A2(n1001), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n704), .A2(n1001), .ZN(n705) );
  XOR2_X1 U796 ( .A(n705), .B(KEYINPUT28), .Z(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U798 ( .A(n708), .B(KEYINPUT29), .ZN(n715) );
  XOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .Z(n709) );
  XNOR2_X1 U800 ( .A(KEYINPUT88), .B(n709), .ZN(n972) );
  NOR2_X1 U801 ( .A1(n972), .A2(n710), .ZN(n713) );
  INV_X1 U802 ( .A(n727), .ZN(n711) );
  XNOR2_X1 U803 ( .A(G1961), .B(KEYINPUT86), .ZN(n961) );
  NOR2_X1 U804 ( .A1(n711), .A2(n961), .ZN(n712) );
  NOR2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n720) );
  NOR2_X1 U806 ( .A1(G301), .A2(n720), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n725) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n727), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n741), .A2(n738), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n716), .A2(G8), .ZN(n717) );
  XNOR2_X1 U811 ( .A(n717), .B(KEYINPUT30), .ZN(n718) );
  NOR2_X1 U812 ( .A1(G168), .A2(n718), .ZN(n719) );
  XNOR2_X1 U813 ( .A(n719), .B(KEYINPUT92), .ZN(n722) );
  AND2_X1 U814 ( .A1(n720), .A2(G301), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U816 ( .A(n723), .B(KEYINPUT31), .ZN(n724) );
  NOR2_X2 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X2 U818 ( .A(n726), .B(KEYINPUT93), .ZN(n739) );
  NAND2_X1 U819 ( .A1(n739), .A2(G286), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n763), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U822 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U823 ( .A(KEYINPUT94), .B(n730), .Z(n731) );
  NOR2_X1 U824 ( .A1(G166), .A2(n731), .ZN(n732) );
  XNOR2_X1 U825 ( .A(n732), .B(KEYINPUT95), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U827 ( .A(n735), .B(KEYINPUT96), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n736), .A2(G8), .ZN(n737) );
  NAND2_X1 U829 ( .A1(G8), .A2(n738), .ZN(n743) );
  INV_X1 U830 ( .A(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n759) );
  NOR2_X1 U834 ( .A1(G2090), .A2(G303), .ZN(n746) );
  XOR2_X1 U835 ( .A(KEYINPUT97), .B(n746), .Z(n747) );
  NAND2_X1 U836 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n759), .A2(n748), .ZN(n749) );
  XNOR2_X1 U838 ( .A(n749), .B(KEYINPUT98), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n750), .A2(n763), .ZN(n754) );
  NOR2_X1 U840 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XOR2_X1 U841 ( .A(n751), .B(KEYINPUT24), .Z(n752) );
  OR2_X1 U842 ( .A1(n763), .A2(n752), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n769) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n1004), .A2(n755), .ZN(n757) );
  INV_X1 U847 ( .A(KEYINPUT33), .ZN(n756) );
  AND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  INV_X1 U851 ( .A(n1002), .ZN(n760) );
  OR2_X1 U852 ( .A1(KEYINPUT33), .A2(n521), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n1004), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n1014) );
  AND2_X1 U858 ( .A1(n767), .A2(n1014), .ZN(n768) );
  INV_X1 U859 ( .A(n771), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n814) );
  XNOR2_X1 U861 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NAND2_X1 U862 ( .A1(G104), .A2(n883), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G140), .A2(n881), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n776), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G128), .A2(n570), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G116), .A2(n878), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n779), .Z(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n782), .ZN(n877) );
  NOR2_X1 U872 ( .A1(n812), .A2(n877), .ZN(n933) );
  NAND2_X1 U873 ( .A1(n814), .A2(n933), .ZN(n810) );
  NAND2_X1 U874 ( .A1(G95), .A2(n883), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G131), .A2(n881), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G119), .A2(n570), .ZN(n786) );
  NAND2_X1 U878 ( .A1(G107), .A2(n878), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n867) );
  INV_X1 U881 ( .A(G1991), .ZN(n968) );
  NOR2_X1 U882 ( .A1(n867), .A2(n968), .ZN(n799) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(KEYINPUT84), .Z(n790) );
  NAND2_X1 U884 ( .A1(G105), .A2(n883), .ZN(n789) );
  XNOR2_X1 U885 ( .A(n790), .B(n789), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G129), .A2(n570), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G117), .A2(n878), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U890 ( .A(KEYINPUT85), .B(n795), .Z(n797) );
  NAND2_X1 U891 ( .A1(n881), .A2(G141), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n863) );
  AND2_X1 U893 ( .A1(n863), .A2(G1996), .ZN(n798) );
  NOR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n916) );
  INV_X1 U895 ( .A(n814), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n916), .A2(n800), .ZN(n807) );
  INV_X1 U897 ( .A(n807), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n810), .A2(n801), .ZN(n802) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n1006) );
  NAND2_X1 U900 ( .A1(n803), .A2(n522), .ZN(n817) );
  NOR2_X1 U901 ( .A1(n863), .A2(G1996), .ZN(n804) );
  XNOR2_X1 U902 ( .A(n804), .B(KEYINPUT100), .ZN(n923) );
  AND2_X1 U903 ( .A1(n968), .A2(n867), .ZN(n930) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U905 ( .A1(n930), .A2(n805), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n923), .A2(n808), .ZN(n809) );
  XNOR2_X1 U908 ( .A(n809), .B(KEYINPUT39), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n812), .A2(n877), .ZN(n915) );
  NAND2_X1 U911 ( .A1(n813), .A2(n915), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n819) );
  XOR2_X1 U914 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n818) );
  XNOR2_X1 U915 ( .A(n819), .B(n818), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U918 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(G188) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XOR2_X1 U925 ( .A(KEYINPUT42), .B(G2090), .Z(n827) );
  XNOR2_X1 U926 ( .A(G2078), .B(G2084), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U928 ( .A(n828), .B(G2100), .Z(n830) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n832) );
  XNOR2_X1 U932 ( .A(KEYINPUT103), .B(G2678), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U934 ( .A(n834), .B(n833), .Z(G227) );
  XNOR2_X1 U935 ( .A(G1991), .B(KEYINPUT41), .ZN(n844) );
  XOR2_X1 U936 ( .A(G1971), .B(G1956), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1961), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U939 ( .A(G1976), .B(G1981), .Z(n838) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1966), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U942 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U943 ( .A(KEYINPUT104), .B(G2474), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G112), .A2(n878), .ZN(n846) );
  NAND2_X1 U947 ( .A1(G136), .A2(n881), .ZN(n845) );
  NAND2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G124), .A2(n570), .ZN(n847) );
  XOR2_X1 U950 ( .A(KEYINPUT44), .B(n847), .Z(n848) );
  XNOR2_X1 U951 ( .A(n848), .B(KEYINPUT105), .ZN(n850) );
  NAND2_X1 U952 ( .A1(G100), .A2(n883), .ZN(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U954 ( .A1(n852), .A2(n851), .ZN(G162) );
  NAND2_X1 U955 ( .A1(n881), .A2(G139), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT110), .ZN(n855) );
  NAND2_X1 U957 ( .A1(G103), .A2(n883), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n570), .A2(G127), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(n856), .Z(n858) );
  NAND2_X1 U961 ( .A1(n878), .A2(G115), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U963 ( .A(KEYINPUT112), .B(n859), .Z(n860) );
  XNOR2_X1 U964 ( .A(KEYINPUT47), .B(n860), .ZN(n861) );
  NOR2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n918) );
  XOR2_X1 U966 ( .A(G160), .B(n863), .Z(n871) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT109), .Z(n865) );
  XNOR2_X1 U968 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n864) );
  XNOR2_X1 U969 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U970 ( .A(n866), .B(KEYINPUT108), .Z(n869) );
  XNOR2_X1 U971 ( .A(n867), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n931), .B(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(G164), .B(G162), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(n918), .B(n875), .Z(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n891) );
  NAND2_X1 U979 ( .A1(G130), .A2(n570), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n889) );
  NAND2_X1 U982 ( .A1(n881), .A2(G142), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n882), .B(KEYINPUT106), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT107), .B(n886), .ZN(n887) );
  XNOR2_X1 U987 ( .A(KEYINPUT45), .B(n887), .ZN(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U990 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U991 ( .A(n893), .B(G286), .Z(n896) );
  XNOR2_X1 U992 ( .A(n894), .B(n998), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n897), .B(G301), .ZN(n898) );
  NOR2_X1 U995 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2438), .B(G2435), .Z(n900) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2430), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(n901), .B(G2454), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2427), .Z(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT102), .B(G2446), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(n907), .B(n906), .Z(n908) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n908), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(n914), .A2(G319), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  INV_X1 U1015 ( .A(n914), .ZN(G401) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n928) );
  XNOR2_X1 U1017 ( .A(G164), .B(G2078), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT115), .ZN(n920) );
  XOR2_X1 U1019 ( .A(G2072), .B(n918), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT50), .B(n921), .ZN(n926) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n936) );
  XOR2_X1 U1027 ( .A(G160), .B(G2084), .Z(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT116), .B(n937), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT52), .B(n938), .Z(n939) );
  XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n990) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n990), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n940), .A2(G29), .ZN(n997) );
  XOR2_X1 U1037 ( .A(G16), .B(KEYINPUT124), .Z(n966) );
  XOR2_X1 U1038 ( .A(G1966), .B(G21), .Z(n952) );
  XNOR2_X1 U1039 ( .A(KEYINPUT125), .B(G1981), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(G6), .ZN(n947) );
  XOR2_X1 U1041 ( .A(KEYINPUT126), .B(G4), .Z(n943) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(n943), .B(n942), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G20), .B(G1956), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n950), .B(KEYINPUT60), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n953), .B(KEYINPUT127), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G1986), .B(G24), .Z(n957) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1057 ( .A(KEYINPUT58), .B(n958), .Z(n959) );
  NAND2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(G5), .B(n961), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n964), .B(KEYINPUT61), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n967), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(G25), .B(n968), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n969), .A2(G28), .ZN(n970) );
  XOR2_X1 U1066 ( .A(KEYINPUT119), .B(n970), .Z(n981) );
  XNOR2_X1 U1067 ( .A(G32), .B(n971), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n972), .B(G27), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G26), .B(G2067), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G33), .B(G2072), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT120), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT53), .B(n982), .Z(n986) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(G34), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n983), .B(KEYINPUT121), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(G2084), .B(n984), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT118), .B(G2090), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(G35), .B(n987), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(n990), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(G29), .A2(n992), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT122), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1024) );
  XOR2_X1 U1089 ( .A(KEYINPUT56), .B(G16), .Z(n1022) );
  XOR2_X1 U1090 ( .A(n998), .B(G1341), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(G171), .B(G1961), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1020) );
  XNOR2_X1 U1093 ( .A(n1001), .B(G1956), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1013) );
  XOR2_X1 U1095 ( .A(n1004), .B(KEYINPUT123), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1007), .B(G1348), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G303), .B(G1971), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G168), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1016), .B(KEYINPUT57), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

