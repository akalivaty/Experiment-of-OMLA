//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n459), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT67), .A3(new_n458), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n465), .B2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n458), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT68), .B1(new_n471), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n459), .A2(new_n481), .A3(new_n458), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n477), .B(new_n479), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n458), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n458), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n459), .A2(KEYINPUT4), .A3(G138), .A4(new_n458), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT69), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n500), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(G50), .A3(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT70), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT7), .Z(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n511), .B2(G89), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n503), .A2(new_n505), .ZN(new_n521));
  INV_X1    g096(.A(new_n501), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n506), .A2(KEYINPUT72), .A3(G63), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n519), .A2(new_n527), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G90), .Z(new_n533));
  NAND3_X1  g108(.A1(new_n506), .A2(new_n510), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n534), .B1(new_n535), .B2(new_n528), .C1(new_n536), .C2(new_n508), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT74), .B(G43), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n529), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n506), .A2(G81), .A3(new_n510), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n542), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT76), .ZN(G188));
  NAND3_X1  g133(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n510), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n506), .A2(G91), .A3(new_n510), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n563), .B(new_n564), .C1(new_n508), .C2(new_n565), .ZN(G299));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n515), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n509), .A2(KEYINPUT77), .A3(new_n512), .A4(new_n514), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G303));
  NAND2_X1  g145(.A1(new_n529), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n506), .A2(G87), .A3(new_n510), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT78), .ZN(G288));
  AND2_X1   g150(.A1(KEYINPUT6), .A2(G651), .ZN(new_n576));
  NOR2_X1   g151(.A1(KEYINPUT6), .A2(G651), .ZN(new_n577));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT79), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n510), .A2(new_n580), .A3(G48), .A4(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n506), .A2(G86), .A3(new_n510), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n506), .B2(G61), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n582), .B(new_n583), .C1(new_n585), .C2(new_n508), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n521), .A2(G61), .A3(new_n522), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n589), .B2(new_n584), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n590), .A2(KEYINPUT80), .A3(new_n583), .A4(new_n582), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n593), .A2(KEYINPUT81), .A3(new_n508), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n511), .A2(G85), .B1(G47), .B2(new_n529), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT81), .B1(new_n593), .B2(new_n508), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n521), .A2(G92), .A3(new_n522), .A4(new_n510), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n506), .A2(new_n601), .A3(G92), .A4(new_n510), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n523), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n598), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n598), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n550), .A2(new_n615), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g199(.A1(new_n480), .A2(new_n482), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n625), .A2(G135), .B1(G123), .B2(new_n476), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT83), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n458), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2438), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2443), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n658), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n666));
  NAND4_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n657), .A4(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n635), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(new_n676), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n678), .A2(new_n680), .A3(new_n683), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n480), .A2(G131), .A3(new_n482), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n476), .A2(G119), .ZN(new_n699));
  OR2_X1    g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n697), .B1(new_n703), .B2(new_n696), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT35), .B(G1991), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n704), .B(new_n705), .Z(new_n706));
  AND2_X1   g281(.A1(KEYINPUT90), .A2(G16), .ZN(new_n707));
  NOR2_X1   g282(.A1(KEYINPUT90), .A2(G16), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(G24), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(G290), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n706), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(G305), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G6), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT32), .B(G1981), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n515), .A2(new_n711), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n709), .A2(G22), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1971), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(G1971), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G1976), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G16), .ZN(new_n735));
  OR2_X1    g310(.A1(G16), .A2(G23), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n574), .B2(new_n719), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT33), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(new_n733), .A3(new_n736), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(KEYINPUT33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n741), .A2(G1976), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n717), .B1(new_n724), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n721), .B(new_n722), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n729), .A2(new_n730), .B1(new_n740), .B2(new_n743), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n747), .A2(KEYINPUT34), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n716), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n696), .A2(G32), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n458), .A2(G105), .A3(G2104), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n754), .B(new_n756), .C1(G129), .C2(new_n476), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n625), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n753), .B1(new_n760), .B2(new_n696), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n630), .A2(G29), .ZN(new_n766));
  OR2_X1    g341(.A1(G5), .A2(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(G1961), .B(new_n767), .C1(G301), .C2(new_n719), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT24), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G34), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n696), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT97), .B(G28), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT30), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n778), .A2(G2084), .B1(new_n696), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n766), .A2(new_n770), .A3(new_n771), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n778), .A2(G2084), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n767), .B1(G301), .B2(new_n719), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n696), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n696), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n786), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n696), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n625), .A2(G140), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n476), .A2(G128), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n696), .ZN(new_n803));
  INV_X1    g378(.A(G2067), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n625), .A2(G139), .ZN(new_n806));
  INV_X1    g381(.A(G127), .ZN(new_n807));
  INV_X1    g382(.A(G115), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n471), .A2(new_n807), .B1(new_n808), .B2(new_n467), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n811), .B1(new_n808), .B2(new_n467), .C1(new_n471), .C2(new_n807), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n810), .A2(G2105), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT25), .Z(new_n815));
  NAND3_X1  g390(.A1(new_n806), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT93), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n806), .A2(new_n813), .A3(new_n818), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G29), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n696), .A2(G33), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT94), .ZN(new_n825));
  INV_X1    g400(.A(G2072), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n821), .A2(new_n827), .A3(new_n823), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n793), .A2(new_n805), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n485), .A2(G29), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT29), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n696), .A2(G35), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g410(.A(G2090), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT23), .B1(new_n709), .B2(G20), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G299), .B2(G16), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n709), .A2(KEYINPUT23), .A3(G20), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n838), .A2(G1956), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(G1956), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n834), .A2(new_n835), .A3(G2090), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n842), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n719), .A2(G4), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n612), .B2(new_n719), .ZN(new_n848));
  INV_X1    g423(.A(G1348), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n762), .A2(new_n764), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n844), .A2(new_n846), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n830), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n825), .A2(new_n828), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT95), .B1(new_n854), .B2(G2072), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n856));
  AOI211_X1 g431(.A(new_n856), .B(new_n826), .C1(new_n825), .C2(new_n828), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n719), .A2(G21), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G168), .B2(new_n719), .ZN(new_n861));
  INV_X1    g436(.A(G1966), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n752), .A2(new_n765), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n709), .A2(G19), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n551), .B2(new_n709), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G1341), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT100), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n746), .A2(new_n749), .ZN(new_n869));
  INV_X1    g444(.A(new_n716), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n751), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI211_X1 g446(.A(KEYINPUT36), .B(new_n716), .C1(new_n746), .C2(new_n749), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n863), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n853), .A2(new_n858), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n877));
  INV_X1    g452(.A(new_n867), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n765), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n879), .ZN(G311));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n878), .A3(new_n765), .ZN(G150));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  INV_X1    g457(.A(G67), .ZN(new_n883));
  AOI211_X1 g458(.A(new_n883), .B(new_n501), .C1(new_n503), .C2(new_n505), .ZN(new_n884));
  NAND2_X1  g459(.A1(G80), .A2(G543), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n882), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(KEYINPUT101), .B(new_n885), .C1(new_n523), .C2(new_n883), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(G651), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n511), .A2(G93), .B1(G55), .B2(new_n529), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n887), .A2(KEYINPUT102), .A3(G651), .A4(new_n888), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G860), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT37), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n551), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n550), .A2(new_n892), .A3(new_n891), .A4(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n611), .A2(new_n619), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n903), .B2(G860), .ZN(G145));
  INV_X1    g479(.A(G142), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT103), .B1(new_n483), .B2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n458), .A2(G118), .ZN(new_n907));
  OAI21_X1  g482(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT104), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n907), .A2(new_n909), .B1(new_n476), .B2(G130), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n480), .A2(new_n911), .A3(new_n482), .A4(G142), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n703), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n702), .A2(new_n906), .A3(new_n910), .A4(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT105), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n633), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n919), .ZN(new_n921));
  INV_X1    g496(.A(new_n633), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n820), .A2(new_n802), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n817), .A2(new_n819), .A3(new_n801), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n495), .A2(new_n496), .A3(new_n489), .A4(new_n488), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n759), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n924), .B2(new_n925), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n920), .B(new_n923), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n925), .ZN(new_n932));
  INV_X1    g507(.A(new_n926), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n759), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n920), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n633), .B1(new_n917), .B2(new_n919), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n935), .B(new_n928), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(G160), .B(new_n485), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n630), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(KEYINPUT106), .A3(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n931), .B2(KEYINPUT107), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n938), .C1(KEYINPUT107), .C2(new_n931), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g525(.A1(new_n894), .A2(G868), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n611), .A2(G299), .ZN(new_n952));
  INV_X1    g527(.A(G299), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(new_n605), .A3(new_n609), .A4(new_n610), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT41), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT41), .B1(new_n952), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n899), .B(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n622), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n899), .B(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n622), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n952), .A2(new_n954), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n967), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT109), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n960), .A2(new_n964), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G290), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n588), .A2(new_n591), .A3(new_n574), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n574), .B1(new_n588), .B2(new_n591), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n515), .B(KEYINPUT110), .Z(new_n979));
  NAND2_X1  g554(.A1(G305), .A2(new_n734), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(G290), .A3(new_n975), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n978), .B2(new_n981), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT42), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n973), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  INV_X1    g562(.A(new_n972), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(new_n965), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(new_n985), .A3(new_n973), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n951), .B1(new_n991), .B2(G868), .ZN(G295));
  AOI21_X1  g567(.A(new_n951), .B1(new_n991), .B2(G868), .ZN(G331));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n515), .B(KEYINPUT110), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n976), .A2(new_n977), .A3(new_n974), .ZN(new_n996));
  AOI21_X1  g571(.A(G290), .B1(new_n980), .B2(new_n975), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G171), .A2(G286), .ZN(new_n1001));
  NAND4_X1  g576(.A1(G301), .A2(new_n530), .A3(new_n527), .A4(new_n519), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n899), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n897), .A2(new_n898), .A3(new_n1003), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n958), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n897), .A2(new_n898), .A3(new_n1003), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n897), .B2(new_n898), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n970), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1000), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n994), .B1(new_n1011), .B2(G37), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT41), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n967), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n955), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1015), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n967), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n984), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G37), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(KEYINPUT112), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1007), .A2(new_n1000), .A3(new_n1010), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1012), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1006), .A2(new_n1005), .B1(new_n971), .B2(new_n969), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n984), .B1(new_n1024), .B2(new_n1016), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1033));
  AND4_X1   g608(.A1(KEYINPUT43), .A2(new_n1025), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT44), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(G397));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n926), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT114), .Z(new_n1039));
  INV_X1    g614(.A(new_n462), .ZN(new_n1040));
  INV_X1    g615(.A(new_n474), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT67), .B1(new_n473), .B2(new_n458), .ZN(new_n1042));
  OAI211_X1 g617(.A(G40), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1039), .A2(KEYINPUT45), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1996), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT115), .A3(new_n760), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n702), .A2(new_n705), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n801), .B(new_n804), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1045), .B2(new_n760), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1044), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1045), .A3(new_n760), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(G2067), .B2(new_n801), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1044), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1046), .A2(KEYINPUT46), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1049), .A2(new_n760), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1044), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1046), .A2(KEYINPUT46), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT47), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1058), .A2(new_n1064), .A3(new_n1061), .A4(new_n1060), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n702), .A2(new_n705), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1044), .B1(new_n1048), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1044), .A2(new_n713), .A3(new_n974), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT48), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1067), .A2(new_n1051), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1057), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT127), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT127), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1057), .A2(new_n1066), .A3(new_n1075), .A4(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT45), .B1(new_n926), .B2(new_n1037), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT120), .B1(new_n1043), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G40), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1080), .B(new_n462), .C1(new_n465), .C2(new_n474), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1078), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1079), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n862), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT50), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1038), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1043), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2084), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n498), .A2(new_n1037), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT116), .B1(new_n1092), .B2(KEYINPUT50), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n1094), .B(new_n1088), .C1(new_n498), .C2(new_n1037), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1090), .B(new_n1091), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1087), .A2(G168), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G168), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(G8), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT51), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1090), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1090), .B(KEYINPUT123), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n784), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT45), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1081), .B1(new_n1108), .B2(new_n1038), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT45), .B1(new_n498), .B2(new_n1037), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1109), .A2(G2078), .A3(new_n1110), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1111), .A2(KEYINPUT53), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1107), .B(new_n1112), .C1(new_n1086), .C2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(G301), .B(KEYINPUT54), .Z(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1100), .A2(new_n1102), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n728), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1103), .B2(G2090), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G8), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n568), .B2(new_n569), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT117), .B(new_n1118), .C1(new_n1103), .C2(G2090), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1121), .A2(new_n1125), .A3(G8), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1123), .B(new_n1124), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1081), .B(new_n1129), .C1(new_n1092), .C2(KEYINPUT50), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1118), .B1(G2090), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G8), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1043), .A2(new_n1038), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(new_n1122), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n574), .A2(new_n732), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT52), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n586), .B(G1981), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1135), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT52), .B1(G288), .B2(new_n732), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(new_n1135), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1140), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1127), .A2(new_n1133), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1039), .A2(KEYINPUT45), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n1150), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(new_n1107), .A3(new_n1115), .A4(new_n1112), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1117), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT122), .B(G2072), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT56), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(G299), .B(KEYINPUT57), .Z(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  INV_X1    g734(.A(G1956), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1130), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1130), .B2(new_n1160), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1157), .B(new_n1158), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1158), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(KEYINPUT124), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT61), .B(new_n1163), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1166), .A2(KEYINPUT126), .A3(new_n1163), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1164), .A2(new_n1173), .A3(new_n1165), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1105), .A2(new_n849), .A3(new_n1106), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1134), .A2(new_n804), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1176), .A2(new_n611), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n611), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT60), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n611), .A2(KEYINPUT60), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT58), .B(G1341), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1134), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1154), .B2(new_n1045), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n551), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n551), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1185), .A2(new_n1190), .B1(KEYINPUT125), .B2(KEYINPUT59), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1181), .A2(new_n1182), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1170), .A2(new_n1175), .A3(new_n1180), .A4(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1163), .B1(new_n1194), .B2(new_n1179), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1153), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1102), .A2(new_n1100), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(KEYINPUT62), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1114), .A2(G171), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1102), .A2(new_n1100), .A3(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1198), .A2(new_n1149), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1127), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1204));
  OR2_X1    g779(.A1(G288), .A2(G1976), .ZN(new_n1205));
  OAI22_X1  g780(.A1(new_n1204), .A2(new_n1205), .B1(G1981), .B2(new_n586), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1203), .A2(new_n1148), .B1(new_n1135), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT63), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1121), .A2(G8), .A3(new_n1126), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1209), .B1(new_n1210), .B2(new_n1128), .ZN(new_n1211));
  AOI211_X1 g786(.A(new_n1122), .B(G286), .C1(new_n1087), .C2(new_n1096), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1211), .A2(new_n1127), .A3(new_n1148), .A4(new_n1212), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1127), .A2(new_n1133), .A3(new_n1148), .A4(new_n1212), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1209), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1196), .A2(new_n1208), .A3(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(G290), .B(G1986), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1044), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1067), .A2(new_n1051), .A3(new_n1069), .A4(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1077), .B1(new_n1217), .B2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g796(.A(new_n673), .B1(new_n651), .B2(new_n652), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n1223), .B1(new_n946), .B2(new_n948), .ZN(new_n1224));
  AND4_X1   g798(.A1(G319), .A2(new_n1030), .A3(new_n694), .A4(new_n1224), .ZN(G308));
  NAND4_X1  g799(.A1(new_n1030), .A2(new_n1224), .A3(G319), .A4(new_n694), .ZN(G225));
endmodule


