

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G651), .A2(G543), .ZN(n652) );
  AND2_X2 U555 ( .A1(n805), .A2(n517), .ZN(n518) );
  NOR2_X2 U556 ( .A1(n698), .A2(n697), .ZN(n700) );
  AND2_X2 U557 ( .A1(n978), .A2(G1348), .ZN(n698) );
  NAND2_X1 U558 ( .A1(n694), .A2(n693), .ZN(n744) );
  NOR2_X1 U559 ( .A1(n813), .A2(n785), .ZN(n805) );
  NOR2_X2 U560 ( .A1(G651), .A2(n535), .ZN(n582) );
  XNOR2_X2 U561 ( .A(KEYINPUT66), .B(n531), .ZN(n583) );
  NOR2_X1 U562 ( .A1(n804), .A2(n519), .ZN(n517) );
  AND2_X1 U563 ( .A1(n803), .A2(n923), .ZN(n519) );
  XNOR2_X1 U564 ( .A(KEYINPUT30), .B(KEYINPUT94), .ZN(n736) );
  XNOR2_X1 U565 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U566 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U567 ( .A1(n734), .A2(n733), .ZN(n753) );
  INV_X1 U568 ( .A(n971), .ZN(n770) );
  NOR2_X1 U569 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U570 ( .A1(G8), .A2(n744), .ZN(n779) );
  NAND2_X1 U571 ( .A1(G160), .A2(G40), .ZN(n692) );
  INV_X1 U572 ( .A(KEYINPUT96), .ZN(n806) );
  NOR2_X2 U573 ( .A1(G2105), .A2(n525), .ZN(n870) );
  XNOR2_X1 U574 ( .A(n521), .B(n520), .ZN(n872) );
  NOR2_X1 U575 ( .A1(n580), .A2(n579), .ZN(n974) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n872), .A2(G137), .ZN(n524) );
  INV_X1 U579 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U580 ( .A1(G101), .A2(n870), .ZN(n522) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n529) );
  AND2_X1 U583 ( .A1(n525), .A2(G2105), .ZN(n866) );
  NAND2_X1 U584 ( .A1(G125), .A2(n866), .ZN(n527) );
  AND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n867) );
  NAND2_X1 U586 ( .A1(G113), .A2(n867), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U588 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U589 ( .A1(n652), .A2(G89), .ZN(n530) );
  XNOR2_X1 U590 ( .A(n530), .B(KEYINPUT4), .ZN(n533) );
  INV_X1 U591 ( .A(G651), .ZN(n536) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n535) );
  NOR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n531) );
  NAND2_X1 U594 ( .A1(G76), .A2(n583), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT5), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G51), .A2(n582), .ZN(n539) );
  NOR2_X1 U598 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n537), .Z(n586) );
  BUF_X1 U600 ( .A(n586), .Z(n651) );
  NAND2_X1 U601 ( .A1(G63), .A2(n651), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n540), .Z(n541) );
  NAND2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U606 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U607 ( .A(G82), .ZN(G220) );
  INV_X1 U608 ( .A(G132), .ZN(G219) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  NOR2_X1 U610 ( .A1(G220), .A2(G219), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT22), .B(n544), .Z(n545) );
  NOR2_X1 U612 ( .A1(G218), .A2(n545), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT81), .B(n546), .Z(n547) );
  NAND2_X1 U614 ( .A1(G96), .A2(n547), .ZN(n915) );
  NAND2_X1 U615 ( .A1(n915), .A2(G2106), .ZN(n552) );
  NAND2_X1 U616 ( .A1(G120), .A2(G69), .ZN(n548) );
  NOR2_X1 U617 ( .A1(G237), .A2(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(KEYINPUT82), .B(n549), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n550), .A2(G108), .ZN(n916) );
  NAND2_X1 U620 ( .A1(n916), .A2(G567), .ZN(n551) );
  AND2_X1 U621 ( .A1(n552), .A2(n551), .ZN(G319) );
  NAND2_X1 U622 ( .A1(G90), .A2(n652), .ZN(n554) );
  NAND2_X1 U623 ( .A1(G77), .A2(n583), .ZN(n553) );
  NAND2_X1 U624 ( .A1(n554), .A2(n553), .ZN(n556) );
  XOR2_X1 U625 ( .A(KEYINPUT68), .B(KEYINPUT9), .Z(n555) );
  XNOR2_X1 U626 ( .A(n556), .B(n555), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G52), .A2(n582), .ZN(n558) );
  NAND2_X1 U628 ( .A1(G64), .A2(n651), .ZN(n557) );
  NAND2_X1 U629 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U630 ( .A(KEYINPUT67), .B(n559), .Z(n560) );
  NOR2_X1 U631 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U632 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U633 ( .A1(G138), .A2(n872), .ZN(n563) );
  NAND2_X1 U634 ( .A1(G102), .A2(n870), .ZN(n562) );
  NAND2_X1 U635 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G126), .A2(n866), .ZN(n565) );
  NAND2_X1 U637 ( .A1(G114), .A2(n867), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U639 ( .A1(n567), .A2(n566), .ZN(G164) );
  XOR2_X1 U640 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n569) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U642 ( .A(n569), .B(n568), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n821) );
  NAND2_X1 U644 ( .A1(n821), .A2(G567), .ZN(n570) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U646 ( .A1(G56), .A2(n651), .ZN(n571) );
  XNOR2_X1 U647 ( .A(n571), .B(KEYINPUT14), .ZN(n574) );
  NAND2_X1 U648 ( .A1(G43), .A2(n582), .ZN(n572) );
  XNOR2_X1 U649 ( .A(n572), .B(KEYINPUT70), .ZN(n573) );
  NAND2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n652), .A2(G81), .ZN(n575) );
  XNOR2_X1 U652 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U653 ( .A1(G68), .A2(n583), .ZN(n576) );
  NAND2_X1 U654 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U655 ( .A(KEYINPUT13), .B(n578), .Z(n579) );
  XNOR2_X1 U656 ( .A(G860), .B(KEYINPUT71), .ZN(n605) );
  INV_X1 U657 ( .A(n605), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n974), .A2(n581), .ZN(G153) );
  XOR2_X1 U659 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  INV_X1 U660 ( .A(G868), .ZN(n668) );
  NOR2_X1 U661 ( .A1(G301), .A2(n668), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G54), .A2(n582), .ZN(n585) );
  NAND2_X1 U663 ( .A1(G79), .A2(n583), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n585), .A2(n584), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G66), .A2(n586), .ZN(n588) );
  NAND2_X1 U666 ( .A1(G92), .A2(n652), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U668 ( .A(n589), .B(KEYINPUT73), .Z(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n592), .Z(n593) );
  XOR2_X2 U671 ( .A(KEYINPUT74), .B(n593), .Z(n978) );
  NOR2_X1 U672 ( .A1(n978), .A2(G868), .ZN(n594) );
  NOR2_X1 U673 ( .A1(n595), .A2(n594), .ZN(G284) );
  XOR2_X1 U674 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U675 ( .A1(G53), .A2(n582), .ZN(n597) );
  NAND2_X1 U676 ( .A1(G65), .A2(n651), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U678 ( .A1(G91), .A2(n652), .ZN(n599) );
  NAND2_X1 U679 ( .A1(G78), .A2(n583), .ZN(n598) );
  NAND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n975) );
  INV_X1 U682 ( .A(n975), .ZN(G299) );
  NOR2_X1 U683 ( .A1(G286), .A2(n668), .ZN(n602) );
  XOR2_X1 U684 ( .A(KEYINPUT75), .B(n602), .Z(n604) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U687 ( .A1(G559), .A2(n605), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n606), .B(KEYINPUT76), .ZN(n607) );
  INV_X1 U689 ( .A(n978), .ZN(n628) );
  NAND2_X1 U690 ( .A1(n607), .A2(n628), .ZN(n608) );
  XNOR2_X1 U691 ( .A(KEYINPUT16), .B(n608), .ZN(G148) );
  NAND2_X1 U692 ( .A1(n974), .A2(n668), .ZN(n609) );
  XNOR2_X1 U693 ( .A(KEYINPUT77), .B(n609), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G868), .A2(n628), .ZN(n610) );
  NOR2_X1 U695 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U696 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U697 ( .A1(n866), .A2(G123), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n613), .B(KEYINPUT18), .ZN(n615) );
  NAND2_X1 U699 ( .A1(G111), .A2(n867), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G135), .A2(n872), .ZN(n617) );
  NAND2_X1 U702 ( .A1(G99), .A2(n870), .ZN(n616) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n922) );
  XNOR2_X1 U705 ( .A(n922), .B(G2096), .ZN(n621) );
  INV_X1 U706 ( .A(G2100), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n621), .A2(n620), .ZN(G156) );
  NAND2_X1 U708 ( .A1(G55), .A2(n582), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G67), .A2(n651), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G93), .A2(n652), .ZN(n625) );
  NAND2_X1 U712 ( .A1(G80), .A2(n583), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n669) );
  NAND2_X1 U715 ( .A1(G559), .A2(n628), .ZN(n666) );
  XOR2_X1 U716 ( .A(n974), .B(n666), .Z(n629) );
  NOR2_X1 U717 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U718 ( .A(n669), .B(n630), .Z(G145) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n631) );
  XNOR2_X1 U720 ( .A(n631), .B(KEYINPUT78), .ZN(n636) );
  NAND2_X1 U721 ( .A1(G49), .A2(n582), .ZN(n633) );
  NAND2_X1 U722 ( .A1(G87), .A2(n535), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U724 ( .A1(n651), .A2(n634), .ZN(n635) );
  NAND2_X1 U725 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G50), .A2(n582), .ZN(n638) );
  NAND2_X1 U727 ( .A1(G62), .A2(n651), .ZN(n637) );
  NAND2_X1 U728 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n652), .A2(G88), .ZN(n639) );
  XOR2_X1 U730 ( .A(KEYINPUT80), .B(n639), .Z(n640) );
  NOR2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U732 ( .A1(G75), .A2(n583), .ZN(n642) );
  NAND2_X1 U733 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  AND2_X1 U735 ( .A1(n652), .A2(G85), .ZN(n647) );
  NAND2_X1 U736 ( .A1(G47), .A2(n582), .ZN(n645) );
  NAND2_X1 U737 ( .A1(G60), .A2(n651), .ZN(n644) );
  NAND2_X1 U738 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U739 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U740 ( .A1(G72), .A2(n583), .ZN(n648) );
  NAND2_X1 U741 ( .A1(n649), .A2(n648), .ZN(G290) );
  NAND2_X1 U742 ( .A1(n583), .A2(G73), .ZN(n650) );
  XOR2_X1 U743 ( .A(KEYINPUT2), .B(n650), .Z(n657) );
  NAND2_X1 U744 ( .A1(G61), .A2(n651), .ZN(n654) );
  NAND2_X1 U745 ( .A1(G86), .A2(n652), .ZN(n653) );
  NAND2_X1 U746 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U747 ( .A(KEYINPUT79), .B(n655), .Z(n656) );
  NOR2_X1 U748 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U749 ( .A1(n582), .A2(G48), .ZN(n658) );
  NAND2_X1 U750 ( .A1(n659), .A2(n658), .ZN(G305) );
  XNOR2_X1 U751 ( .A(G288), .B(KEYINPUT19), .ZN(n661) );
  XNOR2_X1 U752 ( .A(n975), .B(G166), .ZN(n660) );
  XNOR2_X1 U753 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U754 ( .A(n669), .B(n662), .Z(n664) );
  XNOR2_X1 U755 ( .A(G290), .B(n974), .ZN(n663) );
  XNOR2_X1 U756 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U757 ( .A(n665), .B(G305), .Z(n894) );
  XNOR2_X1 U758 ( .A(n666), .B(n894), .ZN(n667) );
  NAND2_X1 U759 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U760 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U761 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U766 ( .A1(n675), .A2(G2072), .ZN(G158) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n676) );
  XNOR2_X1 U768 ( .A(KEYINPUT83), .B(n676), .ZN(n677) );
  NAND2_X1 U769 ( .A1(n677), .A2(G319), .ZN(n678) );
  XOR2_X1 U770 ( .A(KEYINPUT84), .B(n678), .Z(n825) );
  NAND2_X1 U771 ( .A1(G36), .A2(n825), .ZN(G176) );
  NAND2_X1 U772 ( .A1(G128), .A2(n866), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G116), .A2(n867), .ZN(n679) );
  NAND2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U775 ( .A(n681), .B(KEYINPUT35), .ZN(n688) );
  XNOR2_X1 U776 ( .A(KEYINPUT87), .B(KEYINPUT34), .ZN(n686) );
  NAND2_X1 U777 ( .A1(n870), .A2(G104), .ZN(n682) );
  XNOR2_X1 U778 ( .A(n682), .B(KEYINPUT86), .ZN(n684) );
  NAND2_X1 U779 ( .A1(G140), .A2(n872), .ZN(n683) );
  NAND2_X1 U780 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U781 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U783 ( .A(KEYINPUT36), .B(n689), .ZN(n864) );
  XOR2_X1 U784 ( .A(KEYINPUT37), .B(G2067), .Z(n807) );
  NAND2_X1 U785 ( .A1(n864), .A2(n807), .ZN(n937) );
  NOR2_X1 U786 ( .A1(G164), .A2(G1384), .ZN(n694) );
  NOR2_X1 U787 ( .A1(n692), .A2(n694), .ZN(n690) );
  XOR2_X1 U788 ( .A(n690), .B(KEYINPUT85), .Z(n803) );
  INV_X1 U789 ( .A(n803), .ZN(n816) );
  NOR2_X1 U790 ( .A1(n937), .A2(n816), .ZN(n691) );
  XNOR2_X1 U791 ( .A(n691), .B(KEYINPUT88), .ZN(n813) );
  INV_X1 U792 ( .A(n692), .ZN(n693) );
  NOR2_X1 U793 ( .A1(G1981), .A2(G305), .ZN(n695) );
  XOR2_X1 U794 ( .A(n695), .B(KEYINPUT24), .Z(n696) );
  NOR2_X1 U795 ( .A1(n779), .A2(n696), .ZN(n784) );
  INV_X1 U796 ( .A(G1341), .ZN(n998) );
  NOR2_X1 U797 ( .A1(KEYINPUT93), .A2(n998), .ZN(n697) );
  AND2_X1 U798 ( .A1(KEYINPUT26), .A2(n974), .ZN(n699) );
  NAND2_X1 U799 ( .A1(n700), .A2(n699), .ZN(n703) );
  INV_X1 U800 ( .A(n974), .ZN(n701) );
  OR2_X1 U801 ( .A1(n701), .A2(n744), .ZN(n702) );
  AND2_X1 U802 ( .A1(n703), .A2(n702), .ZN(n709) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n978), .ZN(n705) );
  XNOR2_X1 U804 ( .A(G1996), .B(KEYINPUT92), .ZN(n951) );
  NAND2_X1 U805 ( .A1(KEYINPUT26), .A2(n951), .ZN(n704) );
  NAND2_X1 U806 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U807 ( .A1(KEYINPUT93), .A2(n706), .ZN(n707) );
  NOR2_X1 U808 ( .A1(n744), .A2(n707), .ZN(n708) );
  NOR2_X1 U809 ( .A1(n709), .A2(n708), .ZN(n713) );
  OR2_X1 U810 ( .A1(KEYINPUT26), .A2(n951), .ZN(n711) );
  NAND2_X1 U811 ( .A1(KEYINPUT93), .A2(n998), .ZN(n710) );
  AND2_X1 U812 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U813 ( .A1(n713), .A2(n712), .ZN(n723) );
  INV_X1 U814 ( .A(n744), .ZN(n730) );
  NAND2_X1 U815 ( .A1(n730), .A2(G2072), .ZN(n714) );
  XNOR2_X1 U816 ( .A(n714), .B(KEYINPUT27), .ZN(n716) );
  AND2_X1 U817 ( .A1(G1956), .A2(n744), .ZN(n715) );
  NOR2_X1 U818 ( .A1(n716), .A2(n715), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n724), .A2(n975), .ZN(n721) );
  NAND2_X1 U820 ( .A1(G1348), .A2(n744), .ZN(n718) );
  NAND2_X1 U821 ( .A1(G2067), .A2(n730), .ZN(n717) );
  NAND2_X1 U822 ( .A1(n718), .A2(n717), .ZN(n719) );
  OR2_X1 U823 ( .A1(n978), .A2(n719), .ZN(n720) );
  AND2_X1 U824 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U825 ( .A1(n723), .A2(n722), .ZN(n728) );
  NOR2_X1 U826 ( .A1(n724), .A2(n975), .ZN(n726) );
  XNOR2_X1 U827 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n725) );
  XNOR2_X1 U828 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U829 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U830 ( .A(KEYINPUT29), .B(n729), .Z(n734) );
  INV_X1 U831 ( .A(G1961), .ZN(n997) );
  NAND2_X1 U832 ( .A1(n744), .A2(n997), .ZN(n732) );
  XNOR2_X1 U833 ( .A(G2078), .B(KEYINPUT25), .ZN(n950) );
  NAND2_X1 U834 ( .A1(n730), .A2(n950), .ZN(n731) );
  NAND2_X1 U835 ( .A1(n732), .A2(n731), .ZN(n739) );
  NAND2_X1 U836 ( .A1(n739), .A2(G171), .ZN(n733) );
  NOR2_X1 U837 ( .A1(G1966), .A2(n779), .ZN(n754) );
  NOR2_X1 U838 ( .A1(G2084), .A2(n744), .ZN(n756) );
  NOR2_X1 U839 ( .A1(n754), .A2(n756), .ZN(n735) );
  NAND2_X1 U840 ( .A1(G8), .A2(n735), .ZN(n737) );
  NOR2_X1 U841 ( .A1(n738), .A2(G168), .ZN(n741) );
  NOR2_X1 U842 ( .A1(G171), .A2(n739), .ZN(n740) );
  XOR2_X1 U843 ( .A(KEYINPUT31), .B(n742), .Z(n752) );
  NAND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n743) );
  NAND2_X1 U845 ( .A1(n743), .A2(G286), .ZN(n749) );
  NOR2_X1 U846 ( .A1(G1971), .A2(n779), .ZN(n746) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U848 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U849 ( .A1(n747), .A2(G303), .ZN(n748) );
  NAND2_X1 U850 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U851 ( .A1(n750), .A2(G8), .ZN(n751) );
  XNOR2_X1 U852 ( .A(n751), .B(KEYINPUT32), .ZN(n774) );
  AND2_X1 U853 ( .A1(n753), .A2(n752), .ZN(n755) );
  NOR2_X1 U854 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U855 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U856 ( .A1(n758), .A2(n757), .ZN(n775) );
  NAND2_X1 U857 ( .A1(G288), .A2(G1976), .ZN(n759) );
  XOR2_X1 U858 ( .A(KEYINPUT95), .B(n759), .Z(n982) );
  AND2_X1 U859 ( .A1(n775), .A2(n982), .ZN(n760) );
  NAND2_X1 U860 ( .A1(n774), .A2(n760), .ZN(n765) );
  INV_X1 U861 ( .A(n982), .ZN(n762) );
  NOR2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U864 ( .A1(n768), .A2(n761), .ZN(n976) );
  OR2_X1 U865 ( .A1(n762), .A2(n976), .ZN(n763) );
  OR2_X1 U866 ( .A1(n779), .A2(n763), .ZN(n764) );
  NAND2_X1 U867 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U868 ( .A(n766), .B(KEYINPUT64), .ZN(n767) );
  OR2_X2 U869 ( .A1(n767), .A2(KEYINPUT33), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n768), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U871 ( .A1(n769), .A2(n779), .ZN(n771) );
  XOR2_X1 U872 ( .A(G1981), .B(G305), .Z(n971) );
  NAND2_X1 U873 ( .A1(n773), .A2(n772), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n775), .A2(n774), .ZN(n778) );
  NOR2_X1 U875 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U876 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U881 ( .A(G1986), .B(G290), .Z(n983) );
  NOR2_X1 U882 ( .A1(n983), .A2(n816), .ZN(n804) );
  NAND2_X1 U883 ( .A1(G119), .A2(n866), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G131), .A2(n872), .ZN(n787) );
  NAND2_X1 U885 ( .A1(G95), .A2(n870), .ZN(n786) );
  NAND2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U887 ( .A1(G107), .A2(n867), .ZN(n788) );
  XNOR2_X1 U888 ( .A(KEYINPUT89), .B(n788), .ZN(n789) );
  NOR2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U891 ( .A(n793), .B(KEYINPUT90), .ZN(n884) );
  NAND2_X1 U892 ( .A1(n884), .A2(G1991), .ZN(n802) );
  NAND2_X1 U893 ( .A1(G141), .A2(n872), .ZN(n795) );
  NAND2_X1 U894 ( .A1(G129), .A2(n866), .ZN(n794) );
  NAND2_X1 U895 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n870), .A2(G105), .ZN(n796) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(n796), .Z(n797) );
  NOR2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n867), .A2(G117), .ZN(n799) );
  NAND2_X1 U900 ( .A1(n800), .A2(n799), .ZN(n888) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n888), .ZN(n801) );
  NAND2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n923) );
  XNOR2_X1 U903 ( .A(n518), .B(n806), .ZN(n819) );
  NOR2_X1 U904 ( .A1(n864), .A2(n807), .ZN(n928) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n888), .ZN(n919) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n884), .ZN(n924) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U908 ( .A1(n924), .A2(n808), .ZN(n809) );
  NOR2_X1 U909 ( .A1(n519), .A2(n809), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n919), .A2(n810), .ZN(n811) );
  XOR2_X1 U911 ( .A(KEYINPUT39), .B(n811), .Z(n812) );
  NOR2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n928), .A2(n814), .ZN(n815) );
  NOR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT97), .B(n817), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n821), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n822) );
  XNOR2_X1 U920 ( .A(KEYINPUT99), .B(n822), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n823), .A2(G661), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U923 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U924 ( .A(G96), .B(KEYINPUT100), .Z(G221) );
  XOR2_X1 U925 ( .A(KEYINPUT41), .B(G1956), .Z(n827) );
  XNOR2_X1 U926 ( .A(G1986), .B(G1961), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U928 ( .A(n828), .B(KEYINPUT103), .Z(n830) );
  XNOR2_X1 U929 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U931 ( .A(G1976), .B(G1981), .Z(n832) );
  XNOR2_X1 U932 ( .A(G1966), .B(G1971), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U934 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U935 ( .A(KEYINPUT102), .B(G2474), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(G229) );
  XOR2_X1 U937 ( .A(KEYINPUT101), .B(G2090), .Z(n838) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2072), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n839), .B(G2100), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2084), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U943 ( .A(G2096), .B(KEYINPUT43), .Z(n843) );
  XNOR2_X1 U944 ( .A(G2678), .B(KEYINPUT42), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n845), .B(n844), .Z(G227) );
  NAND2_X1 U947 ( .A1(n866), .A2(G124), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U949 ( .A1(G136), .A2(n872), .ZN(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(KEYINPUT104), .B(n849), .Z(n851) );
  NAND2_X1 U952 ( .A1(n867), .A2(G112), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G100), .A2(n870), .ZN(n852) );
  XNOR2_X1 U955 ( .A(KEYINPUT105), .B(n852), .ZN(n853) );
  NOR2_X1 U956 ( .A1(n854), .A2(n853), .ZN(G162) );
  NAND2_X1 U957 ( .A1(n867), .A2(G115), .ZN(n855) );
  XOR2_X1 U958 ( .A(KEYINPUT109), .B(n855), .Z(n857) );
  NAND2_X1 U959 ( .A1(n866), .A2(G127), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT47), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G103), .A2(n870), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n872), .A2(G139), .ZN(n861) );
  XOR2_X1 U965 ( .A(KEYINPUT108), .B(n861), .Z(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n931) );
  XNOR2_X1 U967 ( .A(n864), .B(n931), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(G162), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G130), .A2(n866), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G118), .A2(n867), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n870), .A2(G106), .ZN(n871) );
  XNOR2_X1 U973 ( .A(KEYINPUT106), .B(n871), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n872), .A2(G142), .ZN(n873) );
  XOR2_X1 U975 ( .A(KEYINPUT107), .B(n873), .Z(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n876), .B(KEYINPUT45), .Z(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n890) );
  XOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n882) );
  XNOR2_X1 U981 ( .A(G164), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(n883), .B(n922), .Z(n886) );
  XNOR2_X1 U984 ( .A(G160), .B(n884), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U988 ( .A1(G37), .A2(n891), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n892), .Z(G395) );
  XNOR2_X1 U990 ( .A(G171), .B(n978), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(G286), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G37), .A2(n896), .ZN(n897) );
  XNOR2_X1 U994 ( .A(KEYINPUT112), .B(n897), .ZN(G397) );
  XOR2_X1 U995 ( .A(KEYINPUT98), .B(G2446), .Z(n899) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2454), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n900), .B(G2451), .Z(n902) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1001 ( .A(G2435), .B(G2427), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G2430), .B(G2438), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n907), .ZN(n917) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n917), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1014 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G120), .ZN(G236) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(G325) );
  INV_X1 U1020 ( .A(G325), .ZN(G261) );
  INV_X1 U1021 ( .A(n917), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1029) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1024 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n920), .Z(n930) );
  XOR2_X1 U1026 ( .A(G2084), .B(G160), .Z(n921) );
  NOR2_X1 U1027 ( .A1(n922), .A2(n921), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G2072), .B(n931), .Z(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n932), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G2078), .B(G164), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT117), .B(n933), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(n936), .B(KEYINPUT50), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n944), .A2(G29), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(n945), .ZN(n1027) );
  XOR2_X1 U1045 ( .A(G2067), .B(G26), .Z(n946) );
  NAND2_X1 U1046 ( .A1(G28), .A2(n946), .ZN(n949) );
  XOR2_X1 U1047 ( .A(KEYINPUT121), .B(G2072), .Z(n947) );
  XNOR2_X1 U1048 ( .A(G33), .B(n947), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(n950), .B(G27), .ZN(n953) );
  XOR2_X1 U1051 ( .A(G32), .B(n951), .Z(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(n954), .B(KEYINPUT122), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G25), .B(G1991), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(KEYINPUT120), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n960), .B(KEYINPUT53), .ZN(n963) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1062 ( .A(KEYINPUT119), .B(G2090), .Z(n964) );
  XNOR2_X1 U1063 ( .A(G35), .B(n964), .ZN(n965) );
  NOR2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1065 ( .A(KEYINPUT55), .B(n967), .Z(n968) );
  NOR2_X1 U1066 ( .A1(G29), .A2(n968), .ZN(n969) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(n969), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n970), .A2(G11), .ZN(n1025) );
  XNOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G168), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(KEYINPUT57), .B(n973), .ZN(n994) );
  XNOR2_X1 U1073 ( .A(n974), .B(G1341), .ZN(n991) );
  XNOR2_X1 U1074 ( .A(n975), .B(G1956), .ZN(n977) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n989) );
  XOR2_X1 U1076 ( .A(G171), .B(G1961), .Z(n980) );
  XNOR2_X1 U1077 ( .A(n978), .B(G1348), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(n981), .ZN(n987) );
  AND2_X1 U1080 ( .A1(G303), .A2(G1971), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT125), .B(n992), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1023) );
  INV_X1 U1089 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1090 ( .A(G5), .B(n997), .ZN(n1010) );
  XNOR2_X1 U1091 ( .A(G19), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(G6), .B(G1981), .ZN(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1097 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G21), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(G1986), .B(G24), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1011) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1106 ( .A(G1976), .B(KEYINPUT126), .Z(n1013) );
  XNOR2_X1 U1107 ( .A(G23), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1108 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1109 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(n1029), .B(n1028), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

