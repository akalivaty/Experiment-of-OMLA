

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(n531), .A2(n530), .ZN(G164) );
  XNOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT32), .ZN(n673) );
  XNOR2_X1 U558 ( .A(n674), .B(n673), .ZN(n742) );
  INV_X1 U559 ( .A(KEYINPUT40), .ZN(n775) );
  NOR2_X1 U560 ( .A1(G651), .A2(n586), .ZN(n812) );
  XNOR2_X1 U561 ( .A(n775), .B(KEYINPUT110), .ZN(n776) );
  XNOR2_X1 U562 ( .A(n777), .B(n776), .ZN(G329) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n522), .Z(n893) );
  NAND2_X1 U565 ( .A1(G138), .A2(n893), .ZN(n524) );
  INV_X1 U566 ( .A(G2105), .ZN(n528) );
  AND2_X1 U567 ( .A1(n528), .A2(G2104), .ZN(n892) );
  NAND2_X1 U568 ( .A1(G102), .A2(n892), .ZN(n523) );
  NAND2_X1 U569 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U570 ( .A(KEYINPUT88), .B(n525), .Z(n527) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U572 ( .A1(n898), .A2(G114), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n531) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n528), .ZN(n897) );
  NAND2_X1 U575 ( .A1(G126), .A2(n897), .ZN(n529) );
  XNOR2_X1 U576 ( .A(KEYINPUT87), .B(n529), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G101), .A2(n892), .ZN(n532) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n532), .Z(n535) );
  NAND2_X1 U579 ( .A1(G125), .A2(n897), .ZN(n533) );
  XOR2_X1 U580 ( .A(KEYINPUT65), .B(n533), .Z(n534) );
  NAND2_X1 U581 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U582 ( .A1(n893), .A2(G137), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n898), .A2(G113), .ZN(n536) );
  NAND2_X1 U584 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U585 ( .A1(n539), .A2(n538), .ZN(G160) );
  INV_X1 U586 ( .A(G651), .ZN(n544) );
  NOR2_X1 U587 ( .A1(G543), .A2(n544), .ZN(n540) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n540), .Z(n809) );
  NAND2_X1 U589 ( .A1(G64), .A2(n809), .ZN(n543) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n541) );
  XNOR2_X1 U591 ( .A(KEYINPUT66), .B(n541), .ZN(n586) );
  NAND2_X1 U592 ( .A1(G52), .A2(n812), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n549) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n804) );
  NAND2_X1 U595 ( .A1(G90), .A2(n804), .ZN(n546) );
  NOR2_X1 U596 ( .A1(n544), .A2(n586), .ZN(n805) );
  NAND2_X1 U597 ( .A1(G77), .A2(n805), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U601 ( .A(KEYINPUT68), .B(n550), .Z(G301) );
  INV_X1 U602 ( .A(G301), .ZN(G171) );
  NAND2_X1 U603 ( .A1(G65), .A2(n809), .ZN(n552) );
  NAND2_X1 U604 ( .A1(G78), .A2(n805), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G91), .A2(n804), .ZN(n553) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n553), .ZN(n554) );
  NOR2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n812), .A2(G53), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U611 ( .A1(n804), .A2(G89), .ZN(n558) );
  XNOR2_X1 U612 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U613 ( .A1(G76), .A2(n805), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U615 ( .A(n561), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U616 ( .A1(n812), .A2(G51), .ZN(n562) );
  XNOR2_X1 U617 ( .A(n562), .B(KEYINPUT74), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G63), .A2(n809), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U622 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U623 ( .A1(n812), .A2(G50), .ZN(n570) );
  NAND2_X1 U624 ( .A1(n809), .A2(G62), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U626 ( .A(KEYINPUT83), .B(n571), .ZN(n575) );
  NAND2_X1 U627 ( .A1(G88), .A2(n804), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G75), .A2(n805), .ZN(n572) );
  AND2_X1 U629 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n575), .A2(n574), .ZN(G303) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G60), .A2(n809), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G85), .A2(n804), .ZN(n576) );
  NAND2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U635 ( .A1(G72), .A2(n805), .ZN(n578) );
  XNOR2_X1 U636 ( .A(KEYINPUT67), .B(n578), .ZN(n579) );
  NOR2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n812), .A2(G47), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n582), .A2(n581), .ZN(G290) );
  NAND2_X1 U640 ( .A1(G49), .A2(n812), .ZN(n584) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n583) );
  NAND2_X1 U642 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U643 ( .A1(n809), .A2(n585), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G87), .A2(n586), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n588), .A2(n587), .ZN(G288) );
  NAND2_X1 U646 ( .A1(G61), .A2(n809), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G86), .A2(n804), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U649 ( .A1(n805), .A2(G73), .ZN(n591) );
  XOR2_X1 U650 ( .A(KEYINPUT2), .B(n591), .Z(n592) );
  NOR2_X1 U651 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U652 ( .A(n594), .B(KEYINPUT80), .ZN(n597) );
  NAND2_X1 U653 ( .A1(n812), .A2(G48), .ZN(n595) );
  XOR2_X1 U654 ( .A(KEYINPUT81), .B(n595), .Z(n596) );
  NAND2_X1 U655 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U656 ( .A(n598), .B(KEYINPUT82), .ZN(G305) );
  XOR2_X1 U657 ( .A(G2078), .B(KEYINPUT25), .Z(n959) );
  NOR2_X1 U658 ( .A1(G1384), .A2(G164), .ZN(n600) );
  INV_X1 U659 ( .A(KEYINPUT64), .ZN(n599) );
  XNOR2_X1 U660 ( .A(n600), .B(n599), .ZN(n684) );
  NAND2_X1 U661 ( .A1(G160), .A2(G40), .ZN(n683) );
  OR2_X2 U662 ( .A1(n684), .A2(n683), .ZN(n661) );
  XOR2_X1 U663 ( .A(n661), .B(KEYINPUT98), .Z(n613) );
  INV_X1 U664 ( .A(n613), .ZN(n605) );
  NOR2_X1 U665 ( .A1(n959), .A2(n605), .ZN(n603) );
  NOR2_X1 U666 ( .A1(n683), .A2(n684), .ZN(n601) );
  XOR2_X1 U667 ( .A(G1961), .B(KEYINPUT97), .Z(n1008) );
  NOR2_X1 U668 ( .A1(n601), .A2(n1008), .ZN(n602) );
  NOR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT99), .B(n604), .ZN(n656) );
  NAND2_X1 U671 ( .A1(n656), .A2(G171), .ZN(n651) );
  INV_X1 U672 ( .A(G299), .ZN(n985) );
  NAND2_X1 U673 ( .A1(n605), .A2(G1956), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n606), .B(KEYINPUT100), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G2072), .A2(n613), .ZN(n607) );
  XOR2_X1 U676 ( .A(KEYINPUT27), .B(n607), .Z(n608) );
  NAND2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n610), .B(KEYINPUT101), .ZN(n612) );
  NOR2_X1 U679 ( .A1(n985), .A2(n612), .ZN(n611) );
  XOR2_X1 U680 ( .A(n611), .B(KEYINPUT28), .Z(n648) );
  NAND2_X1 U681 ( .A1(n985), .A2(n612), .ZN(n646) );
  NAND2_X1 U682 ( .A1(n613), .A2(G2067), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G1348), .A2(n661), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n640) );
  XOR2_X1 U685 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n617) );
  NAND2_X1 U686 ( .A1(G56), .A2(n809), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n804), .A2(G81), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT12), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G68), .A2(n805), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U692 ( .A(KEYINPUT13), .B(n621), .Z(n622) );
  NOR2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n812), .A2(G43), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n988) );
  XOR2_X1 U696 ( .A(G1996), .B(KEYINPUT102), .Z(n958) );
  NOR2_X1 U697 ( .A1(n661), .A2(n958), .ZN(n626) );
  XOR2_X1 U698 ( .A(n626), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U699 ( .A1(n661), .A2(G1341), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n988), .A2(n629), .ZN(n642) );
  NAND2_X1 U702 ( .A1(G66), .A2(n809), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G92), .A2(n804), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U705 ( .A1(G54), .A2(n812), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G79), .A2(n805), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U709 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n637), .B(n636), .ZN(n638) );
  XOR2_X1 U711 ( .A(KEYINPUT15), .B(n638), .Z(n908) );
  INV_X1 U712 ( .A(n908), .ZN(n989) );
  NAND2_X1 U713 ( .A1(n642), .A2(n989), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U715 ( .A(KEYINPUT103), .B(n641), .Z(n644) );
  OR2_X1 U716 ( .A1(n989), .A2(n642), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U720 ( .A(n649), .B(KEYINPUT29), .Z(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n680) );
  NAND2_X1 U722 ( .A1(G8), .A2(n661), .ZN(n758) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n758), .ZN(n678) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n661), .ZN(n675) );
  NOR2_X1 U725 ( .A1(n678), .A2(n675), .ZN(n652) );
  XNOR2_X1 U726 ( .A(KEYINPUT104), .B(n652), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n653), .A2(G8), .ZN(n654) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n654), .ZN(n655) );
  NOR2_X1 U729 ( .A1(G168), .A2(n655), .ZN(n658) );
  NOR2_X1 U730 ( .A1(G171), .A2(n656), .ZN(n657) );
  NOR2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT31), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT105), .ZN(n679) );
  INV_X1 U734 ( .A(G8), .ZN(n666) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n758), .ZN(n663) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n661), .ZN(n662) );
  NOR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n664), .A2(G303), .ZN(n665) );
  OR2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n668) );
  AND2_X1 U740 ( .A1(n679), .A2(n668), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n680), .A2(n667), .ZN(n672) );
  INV_X1 U742 ( .A(n668), .ZN(n670) );
  AND2_X1 U743 ( .A1(G286), .A2(G8), .ZN(n669) );
  OR2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U746 ( .A1(G8), .A2(n675), .ZN(n676) );
  XOR2_X1 U747 ( .A(KEYINPUT96), .B(n676), .Z(n677) );
  NOR2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n738) );
  INV_X1 U751 ( .A(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n705) );
  INV_X1 U753 ( .A(n705), .ZN(n768) );
  NAND2_X1 U754 ( .A1(G105), .A2(n892), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT94), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n687), .B(KEYINPUT38), .ZN(n689) );
  NAND2_X1 U757 ( .A1(G141), .A2(n893), .ZN(n688) );
  NAND2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U759 ( .A1(G129), .A2(n897), .ZN(n690) );
  XNOR2_X1 U760 ( .A(KEYINPUT93), .B(n690), .ZN(n691) );
  NOR2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n898), .A2(G117), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n885) );
  NOR2_X1 U764 ( .A1(G1996), .A2(n885), .ZN(n938) );
  NAND2_X1 U765 ( .A1(G1996), .A2(n885), .ZN(n695) );
  XNOR2_X1 U766 ( .A(n695), .B(KEYINPUT95), .ZN(n704) );
  NAND2_X1 U767 ( .A1(G95), .A2(n892), .ZN(n697) );
  NAND2_X1 U768 ( .A1(G131), .A2(n893), .ZN(n696) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U770 ( .A(KEYINPUT92), .B(n698), .Z(n702) );
  NAND2_X1 U771 ( .A1(G119), .A2(n897), .ZN(n700) );
  NAND2_X1 U772 ( .A1(G107), .A2(n898), .ZN(n699) );
  AND2_X1 U773 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U774 ( .A1(n702), .A2(n701), .ZN(n889) );
  AND2_X1 U775 ( .A1(G1991), .A2(n889), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n948) );
  NOR2_X1 U777 ( .A1(n948), .A2(n705), .ZN(n765) );
  NOR2_X1 U778 ( .A1(G1986), .A2(G290), .ZN(n706) );
  NOR2_X1 U779 ( .A1(G1991), .A2(n889), .ZN(n946) );
  NOR2_X1 U780 ( .A1(n706), .A2(n946), .ZN(n707) );
  NOR2_X1 U781 ( .A1(n765), .A2(n707), .ZN(n708) );
  NOR2_X1 U782 ( .A1(n938), .A2(n708), .ZN(n709) );
  XNOR2_X1 U783 ( .A(n709), .B(KEYINPUT39), .ZN(n722) );
  NAND2_X1 U784 ( .A1(n892), .A2(G104), .ZN(n710) );
  XOR2_X1 U785 ( .A(KEYINPUT89), .B(n710), .Z(n712) );
  NAND2_X1 U786 ( .A1(n893), .A2(G140), .ZN(n711) );
  NAND2_X1 U787 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U788 ( .A(KEYINPUT34), .B(n713), .ZN(n718) );
  NAND2_X1 U789 ( .A1(G128), .A2(n897), .ZN(n715) );
  NAND2_X1 U790 ( .A1(G116), .A2(n898), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U792 ( .A(n716), .B(KEYINPUT35), .Z(n717) );
  NOR2_X1 U793 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U794 ( .A(KEYINPUT36), .B(n719), .Z(n720) );
  XOR2_X1 U795 ( .A(KEYINPUT90), .B(n720), .Z(n884) );
  XNOR2_X1 U796 ( .A(KEYINPUT37), .B(G2067), .ZN(n723) );
  OR2_X1 U797 ( .A1(n884), .A2(n723), .ZN(n721) );
  XNOR2_X1 U798 ( .A(n721), .B(KEYINPUT91), .ZN(n950) );
  NAND2_X1 U799 ( .A1(n768), .A2(n950), .ZN(n766) );
  NAND2_X1 U800 ( .A1(n722), .A2(n766), .ZN(n724) );
  NAND2_X1 U801 ( .A1(n884), .A2(n723), .ZN(n954) );
  NAND2_X1 U802 ( .A1(n724), .A2(n954), .ZN(n725) );
  NAND2_X1 U803 ( .A1(n768), .A2(n725), .ZN(n726) );
  XNOR2_X1 U804 ( .A(n726), .B(KEYINPUT109), .ZN(n772) );
  OR2_X1 U805 ( .A1(n772), .A2(n758), .ZN(n728) );
  AND2_X1 U806 ( .A1(n738), .A2(n728), .ZN(n727) );
  NAND2_X1 U807 ( .A1(n742), .A2(n727), .ZN(n735) );
  INV_X1 U808 ( .A(n728), .ZN(n733) );
  NOR2_X1 U809 ( .A1(G2090), .A2(G303), .ZN(n729) );
  NAND2_X1 U810 ( .A1(G8), .A2(n729), .ZN(n731) );
  INV_X1 U811 ( .A(n772), .ZN(n730) );
  AND2_X1 U812 ( .A1(n731), .A2(n730), .ZN(n732) );
  OR2_X1 U813 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U814 ( .A1(n735), .A2(n734), .ZN(n764) );
  NAND2_X1 U815 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U816 ( .A(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n745) );
  INV_X1 U818 ( .A(n745), .ZN(n994) );
  OR2_X1 U819 ( .A1(n758), .A2(n994), .ZN(n736) );
  NOR2_X1 U820 ( .A1(n751), .A2(n736), .ZN(n737) );
  XOR2_X1 U821 ( .A(n737), .B(KEYINPUT108), .Z(n750) );
  AND2_X1 U822 ( .A1(n995), .A2(n750), .ZN(n743) );
  AND2_X1 U823 ( .A1(n738), .A2(n743), .ZN(n740) );
  XNOR2_X1 U824 ( .A(G1981), .B(G305), .ZN(n983) );
  INV_X1 U825 ( .A(n983), .ZN(n739) );
  AND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n762) );
  INV_X1 U828 ( .A(n743), .ZN(n749) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n744) );
  XOR2_X1 U830 ( .A(KEYINPUT107), .B(n744), .Z(n746) );
  NOR2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U832 ( .A1(n758), .A2(n747), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n754) );
  INV_X1 U834 ( .A(n750), .ZN(n752) );
  NOR2_X1 U835 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U836 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U837 ( .A1(n983), .A2(n755), .ZN(n760) );
  NOR2_X1 U838 ( .A1(G1981), .A2(G305), .ZN(n756) );
  XOR2_X1 U839 ( .A(n756), .B(KEYINPUT24), .Z(n757) );
  NOR2_X1 U840 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U841 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U842 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U843 ( .A1(n764), .A2(n763), .ZN(n774) );
  INV_X1 U844 ( .A(n765), .ZN(n767) );
  AND2_X1 U845 ( .A1(n767), .A2(n766), .ZN(n770) );
  XNOR2_X1 U846 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U847 ( .A1(n768), .A2(n987), .ZN(n769) );
  AND2_X1 U848 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U849 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U850 ( .A1(n774), .A2(n773), .ZN(n777) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U852 ( .A(G57), .ZN(G237) );
  INV_X1 U853 ( .A(G132), .ZN(G219) );
  INV_X1 U854 ( .A(G82), .ZN(G220) );
  NAND2_X1 U855 ( .A1(G7), .A2(G661), .ZN(n778) );
  XOR2_X1 U856 ( .A(n778), .B(KEYINPUT10), .Z(n842) );
  NAND2_X1 U857 ( .A1(n842), .A2(G567), .ZN(n779) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n803) );
  OR2_X1 U860 ( .A1(n988), .A2(n803), .ZN(G153) );
  INV_X1 U861 ( .A(G868), .ZN(n783) );
  NOR2_X1 U862 ( .A1(n783), .A2(G171), .ZN(n780) );
  XNOR2_X1 U863 ( .A(n780), .B(KEYINPUT71), .ZN(n782) );
  NAND2_X1 U864 ( .A1(n783), .A2(n908), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n782), .A2(n781), .ZN(G284) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U867 ( .A1(G286), .A2(n783), .ZN(n784) );
  NOR2_X1 U868 ( .A1(n785), .A2(n784), .ZN(G297) );
  NAND2_X1 U869 ( .A1(n803), .A2(G559), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n786), .A2(n989), .ZN(n787) );
  XNOR2_X1 U871 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U872 ( .A1(G868), .A2(n988), .ZN(n790) );
  NAND2_X1 U873 ( .A1(n989), .A2(G868), .ZN(n788) );
  NOR2_X1 U874 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n897), .ZN(n791) );
  XNOR2_X1 U877 ( .A(n791), .B(KEYINPUT18), .ZN(n799) );
  NAND2_X1 U878 ( .A1(n892), .A2(G99), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n792), .B(KEYINPUT76), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G111), .A2(n898), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G135), .A2(n893), .ZN(n795) );
  XNOR2_X1 U883 ( .A(KEYINPUT75), .B(n795), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n943) );
  XNOR2_X1 U886 ( .A(G2096), .B(n943), .ZN(n800) );
  NOR2_X1 U887 ( .A1(n800), .A2(G2100), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n801), .B(KEYINPUT77), .ZN(G156) );
  NAND2_X1 U889 ( .A1(n989), .A2(G559), .ZN(n802) );
  XOR2_X1 U890 ( .A(n988), .B(n802), .Z(n824) );
  NAND2_X1 U891 ( .A1(n803), .A2(n824), .ZN(n816) );
  NAND2_X1 U892 ( .A1(G93), .A2(n804), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G80), .A2(n805), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U895 ( .A(KEYINPUT78), .B(n808), .Z(n811) );
  NAND2_X1 U896 ( .A1(n809), .A2(G67), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G55), .A2(n812), .ZN(n813) );
  XNOR2_X1 U899 ( .A(KEYINPUT79), .B(n813), .ZN(n814) );
  NOR2_X1 U900 ( .A1(n815), .A2(n814), .ZN(n826) );
  XOR2_X1 U901 ( .A(n816), .B(n826), .Z(G145) );
  XNOR2_X1 U902 ( .A(G305), .B(n826), .ZN(n823) );
  XNOR2_X1 U903 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n818) );
  XNOR2_X1 U904 ( .A(G288), .B(KEYINPUT19), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n818), .B(n817), .ZN(n819) );
  XNOR2_X1 U906 ( .A(G290), .B(n819), .ZN(n821) );
  XOR2_X1 U907 ( .A(G303), .B(n985), .Z(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n823), .B(n822), .ZN(n907) );
  XNOR2_X1 U910 ( .A(n824), .B(n907), .ZN(n825) );
  NAND2_X1 U911 ( .A1(n825), .A2(G868), .ZN(n828) );
  OR2_X1 U912 ( .A1(G868), .A2(n826), .ZN(n827) );
  NAND2_X1 U913 ( .A1(n828), .A2(n827), .ZN(G295) );
  NAND2_X1 U914 ( .A1(G2078), .A2(G2084), .ZN(n829) );
  XOR2_X1 U915 ( .A(KEYINPUT20), .B(n829), .Z(n830) );
  NAND2_X1 U916 ( .A1(G2090), .A2(n830), .ZN(n832) );
  XNOR2_X1 U917 ( .A(KEYINPUT86), .B(KEYINPUT21), .ZN(n831) );
  XNOR2_X1 U918 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U919 ( .A1(G2072), .A2(n833), .ZN(G158) );
  XNOR2_X1 U920 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U921 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U922 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U923 ( .A1(G218), .A2(n835), .ZN(n836) );
  NAND2_X1 U924 ( .A1(G96), .A2(n836), .ZN(n929) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n929), .ZN(n840) );
  NAND2_X1 U926 ( .A1(G69), .A2(G120), .ZN(n837) );
  NOR2_X1 U927 ( .A1(G237), .A2(n837), .ZN(n838) );
  NAND2_X1 U928 ( .A1(G108), .A2(n838), .ZN(n930) );
  NAND2_X1 U929 ( .A1(G567), .A2(n930), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n863) );
  NAND2_X1 U931 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n863), .A2(n841), .ZN(n845) );
  NAND2_X1 U933 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n842), .ZN(G217) );
  INV_X1 U935 ( .A(n842), .ZN(G223) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(G188) );
  XOR2_X1 U940 ( .A(G1986), .B(G1981), .Z(n847) );
  XNOR2_X1 U941 ( .A(G1956), .B(G1966), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U943 ( .A(n848), .B(G2474), .Z(n850) );
  XNOR2_X1 U944 ( .A(G1991), .B(G1996), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1976), .Z(n852) );
  XNOR2_X1 U947 ( .A(G1971), .B(G1961), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U949 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U950 ( .A(G2100), .B(G2096), .Z(n856) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2072), .Z(n858) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2090), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U956 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(G227) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(n863), .ZN(G319) );
  NAND2_X1 U960 ( .A1(G124), .A2(n897), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U962 ( .A1(n892), .A2(G100), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U964 ( .A1(G136), .A2(n893), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G112), .A2(n898), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U967 ( .A1(n870), .A2(n869), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n872) );
  XNOR2_X1 U969 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT48), .B(n873), .Z(n883) );
  NAND2_X1 U972 ( .A1(G130), .A2(n897), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G118), .A2(n898), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U975 ( .A1(G106), .A2(n892), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G142), .A2(n893), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(n878), .B(KEYINPUT45), .Z(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(n943), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U984 ( .A(n888), .B(G162), .Z(n891) );
  XOR2_X1 U985 ( .A(n889), .B(G160), .Z(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n905) );
  NAND2_X1 U987 ( .A1(G103), .A2(n892), .ZN(n895) );
  NAND2_X1 U988 ( .A1(G139), .A2(n893), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(KEYINPUT113), .B(n896), .Z(n903) );
  NAND2_X1 U991 ( .A1(G127), .A2(n897), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U993 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U995 ( .A1(n903), .A2(n902), .ZN(n932) );
  XNOR2_X1 U996 ( .A(n932), .B(G164), .ZN(n904) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U998 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n988), .B(n907), .ZN(n910) );
  XOR2_X1 U1000 ( .A(G171), .B(n908), .Z(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1002 ( .A(n911), .B(G286), .ZN(n912) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1004 ( .A(KEYINPUT116), .B(n913), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1006 ( .A(n914), .B(KEYINPUT49), .ZN(n926) );
  XOR2_X1 U1007 ( .A(G2451), .B(G2430), .Z(n916) );
  XNOR2_X1 U1008 ( .A(G2438), .B(G2443), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n916), .B(n915), .ZN(n922) );
  XOR2_X1 U1010 ( .A(G2435), .B(G2454), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1013 ( .A(G2446), .B(G2427), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1015 ( .A(n922), .B(n921), .Z(n923) );
  NAND2_X1 U1016 ( .A1(G14), .A2(n923), .ZN(n931) );
  NAND2_X1 U1017 ( .A1(n931), .A2(G319), .ZN(n924) );
  XOR2_X1 U1018 ( .A(KEYINPUT117), .B(n924), .Z(n925) );
  NOR2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(G225) );
  XOR2_X1 U1022 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1024 ( .A(G120), .ZN(G236) );
  INV_X1 U1025 ( .A(G96), .ZN(G221) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(G325) );
  INV_X1 U1028 ( .A(G325), .ZN(G261) );
  INV_X1 U1029 ( .A(G303), .ZN(G166) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  INV_X1 U1031 ( .A(n931), .ZN(G401) );
  XNOR2_X1 U1032 ( .A(G2072), .B(n932), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n933), .B(KEYINPUT121), .ZN(n935) );
  XOR2_X1 U1034 ( .A(G2078), .B(G164), .Z(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT50), .B(n936), .ZN(n942) );
  XOR2_X1 U1037 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT120), .B(n940), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(G160), .B(G2084), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT119), .B(n951), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n956), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n957), .A2(G29), .ZN(n1036) );
  XOR2_X1 U1052 ( .A(n958), .B(G32), .Z(n961) );
  XNOR2_X1 U1053 ( .A(n959), .B(G27), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n971) );
  XOR2_X1 U1055 ( .A(G25), .B(G1991), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(G28), .ZN(n969) );
  XOR2_X1 U1057 ( .A(G2072), .B(KEYINPUT123), .Z(n963) );
  XNOR2_X1 U1058 ( .A(G33), .B(n963), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT122), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1062 ( .A(KEYINPUT124), .B(n967), .Z(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT53), .ZN(n975) );
  XOR2_X1 U1066 ( .A(G2084), .B(G34), .Z(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT54), .B(n973), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G35), .B(G2090), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1071 ( .A(KEYINPUT125), .B(n978), .Z(n979) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n979), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(KEYINPUT55), .B(n980), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(G11), .ZN(n1034) );
  INV_X1 U1075 ( .A(G16), .ZN(n1030) );
  XOR2_X1 U1076 ( .A(n1030), .B(KEYINPUT56), .Z(n1007) );
  XOR2_X1 U1077 ( .A(G1966), .B(G168), .Z(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n984), .Z(n1005) );
  XOR2_X1 U1080 ( .A(G1961), .B(G301), .Z(n1000) );
  XOR2_X1 U1081 ( .A(G1956), .B(n985), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n988), .B(G1341), .ZN(n991) );
  XOR2_X1 U1084 ( .A(n989), .B(G1348), .Z(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT126), .B(n996), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G166), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT127), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1032) );
  XNOR2_X1 U1096 ( .A(n1008), .B(G5), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G21), .B(G1966), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1020) );
  XOR2_X1 U1099 ( .A(G1348), .B(KEYINPUT59), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G20), .B(G1956), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G1341), .B(G19), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G1981), .B(G6), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1018), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(G1971), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1112 ( .A(G1986), .B(G24), .Z(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1037), .ZN(G150) );
  INV_X1 U1122 ( .A(G150), .ZN(G311) );
endmodule

