//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT82), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n187), .A2(new_n188), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(KEYINPUT84), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n193));
  INV_X1    g007(.A(G110), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G122), .ZN(new_n195));
  INV_X1    g009(.A(G122), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G110), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT82), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n189), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n192), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n192), .B2(new_n199), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G116), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G113), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(G119), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n212), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n211), .A2(new_n218), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n224), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(G104), .ZN(new_n228));
  INV_X1    g042(.A(G101), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(G107), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n225), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n224), .A2(G107), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n227), .A2(G104), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n223), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G143), .ZN(new_n238));
  INV_X1    g052(.A(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n241), .A2(KEYINPUT1), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  AOI21_X1  g058(.A(G128), .B1(new_n238), .B2(new_n240), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n239), .A2(KEYINPUT1), .A3(G146), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G143), .B(G146), .ZN(new_n249));
  OAI211_X1 g063(.A(KEYINPUT66), .B(new_n246), .C1(new_n249), .C2(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n243), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n241), .A2(new_n258), .A3(KEYINPUT64), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G224), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT7), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n203), .A2(new_n236), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n253), .A2(new_n261), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT85), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT7), .A4(new_n264), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n225), .A2(new_n228), .A3(new_n230), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G101), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n270), .A2(KEYINPUT79), .A3(new_n271), .A4(G101), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n211), .A2(new_n218), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n209), .A2(new_n210), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(G101), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n219), .A2(new_n222), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n231), .A2(new_n234), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT81), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n190), .A2(new_n191), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n223), .A2(new_n288), .A3(new_n235), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n282), .A2(new_n286), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n261), .A4(new_n264), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n266), .A2(new_n269), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n286), .A3(new_n289), .ZN(new_n296));
  INV_X1    g110(.A(new_n287), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT6), .A4(new_n290), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n290), .A2(KEYINPUT6), .ZN(new_n301));
  AND4_X1   g115(.A1(new_n288), .A2(new_n277), .A3(new_n235), .A4(new_n283), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n288), .B1(new_n223), .B2(new_n235), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n304), .B2(new_n282), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT6), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n296), .A2(new_n307), .A3(new_n297), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT83), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n300), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n262), .B(new_n264), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n295), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G210), .B1(G237), .B2(G902), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT87), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n313), .B2(KEYINPUT86), .ZN(new_n317));
  OAI211_X1 g131(.A(KEYINPUT83), .B(new_n308), .C1(new_n301), .C2(new_n305), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n311), .B1(new_n318), .B2(new_n300), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(new_n320), .A3(new_n295), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n315), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n320), .B1(new_n319), .B2(new_n295), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(KEYINPUT87), .A3(new_n316), .A4(new_n325), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n322), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n249), .A2(new_n328), .A3(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n241), .A2(new_n242), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT66), .B1(new_n330), .B2(new_n246), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n245), .A2(new_n244), .A3(new_n247), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT10), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n285), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n330), .A3(new_n246), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n235), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n333), .A2(new_n335), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT11), .ZN(new_n340));
  INV_X1    g154(.A(G134), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n339), .B(new_n340), .C1(new_n341), .C2(G137), .ZN(new_n342));
  INV_X1    g156(.A(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT11), .A3(G134), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(G137), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(G134), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n339), .B1(new_n347), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g162(.A(G131), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n344), .A2(new_n345), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n340), .B1(new_n341), .B2(G137), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT65), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .A4(new_n342), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n256), .A2(new_n259), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n276), .A2(new_n356), .A3(new_n281), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n338), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n329), .B(new_n285), .C1(new_n331), .C2(new_n332), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n337), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n349), .A2(new_n354), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n360), .A2(KEYINPUT12), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT12), .B1(new_n360), .B2(new_n361), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n263), .A2(G227), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n338), .A2(new_n357), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n361), .ZN(new_n370));
  INV_X1    g184(.A(new_n367), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n358), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n294), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G469), .ZN(new_n375));
  INV_X1    g189(.A(new_n358), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n355), .B1(new_n338), .B2(new_n357), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n367), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n358), .B(new_n371), .C1(new_n362), .C2(new_n363), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n381));
  INV_X1    g195(.A(G469), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n375), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  OAI21_X1  g200(.A(G221), .B1(new_n386), .B2(G902), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n263), .A2(G952), .ZN(new_n389));
  INV_X1    g203(.A(G234), .ZN(new_n390));
  INV_X1    g204(.A(G237), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n294), .B(new_n263), .C1(G234), .C2(G237), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n386), .A2(new_n397), .A3(G953), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT94), .B1(new_n196), .B2(G116), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT94), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n207), .A3(G122), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n402), .A2(KEYINPUT14), .B1(G116), .B2(new_n196), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(KEYINPUT96), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(KEYINPUT96), .B2(new_n404), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n239), .A2(G128), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT95), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n239), .A2(G128), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n410), .A2(G134), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n408), .B(KEYINPUT95), .ZN(new_n413));
  INV_X1    g227(.A(new_n411), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n341), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n402), .B1(new_n207), .B2(G122), .ZN(new_n416));
  OAI22_X1  g230(.A1(new_n412), .A2(new_n415), .B1(G107), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n341), .A3(new_n414), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n416), .A2(G107), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n416), .A2(G107), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT13), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n411), .B1(new_n413), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n341), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n398), .B1(new_n419), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n417), .B1(new_n406), .B2(G107), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n423), .A2(new_n427), .ZN(new_n431));
  INV_X1    g245(.A(new_n398), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n294), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n419), .A2(new_n428), .A3(new_n398), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n432), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n440), .B(new_n294), .C1(KEYINPUT15), .C2(new_n435), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G113), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n224), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n391), .A2(new_n263), .A3(G214), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n239), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n391), .A2(new_n263), .A3(G143), .A4(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT88), .ZN(new_n449));
  AND2_X1   g263(.A1(KEYINPUT18), .A2(G131), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G125), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n252), .A2(G140), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n237), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT76), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT76), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .A4(new_n237), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(KEYINPUT72), .A2(G125), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT73), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G140), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT73), .B1(new_n452), .B2(G125), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n452), .A2(KEYINPUT72), .A3(G125), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n451), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT16), .B1(new_n452), .B2(G125), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n465), .B2(KEYINPUT16), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G146), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT93), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(KEYINPUT16), .ZN(new_n473));
  INV_X1    g287(.A(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n237), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n448), .A2(KEYINPUT90), .A3(G131), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT90), .B1(new_n448), .B2(G131), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT17), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n448), .A2(G131), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT89), .B1(new_n448), .B2(G131), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n446), .A2(new_n490), .A3(new_n351), .A4(new_n447), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n488), .A2(new_n482), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n485), .B1(new_n492), .B2(KEYINPUT17), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n444), .B(new_n468), .C1(new_n481), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n483), .A2(new_n484), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n489), .A4(new_n491), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n498), .A2(new_n472), .A3(new_n480), .A4(new_n485), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n444), .B1(new_n499), .B2(new_n468), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n294), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G475), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n465), .A2(KEYINPUT19), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT19), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n453), .A2(new_n454), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n504), .A2(new_n237), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n237), .B1(new_n473), .B2(new_n474), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT91), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n237), .A3(new_n506), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n511), .C1(new_n237), .C2(new_n470), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n492), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT92), .A3(new_n468), .ZN(new_n514));
  INV_X1    g328(.A(new_n444), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT92), .B1(new_n513), .B2(new_n468), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n494), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n503), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n518), .A2(new_n503), .A3(new_n519), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n442), .B(new_n502), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n388), .A2(new_n396), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n327), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G472), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n347), .A2(new_n345), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G131), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n354), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n251), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n260), .B1(new_n354), .B2(new_n349), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n279), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n361), .A2(new_n356), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n277), .A2(new_n278), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n534), .C1(new_n251), .C2(new_n529), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n526), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n535), .A2(new_n526), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G210), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n540), .A2(G237), .A3(G953), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n537), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT30), .B1(new_n530), .B2(new_n531), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n533), .B(new_n549), .C1(new_n251), .C2(new_n529), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n534), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n535), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n546), .B(new_n547), .C1(new_n553), .C2(new_n545), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n536), .A2(new_n538), .A3(new_n544), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n555), .B2(KEYINPUT29), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n525), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR4_X1   g371(.A1(new_n551), .A2(KEYINPUT31), .A3(new_n552), .A4(new_n544), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n544), .B1(new_n536), .B2(new_n538), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n545), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT32), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT32), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n559), .A2(new_n560), .B1(new_n553), .B2(new_n545), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n567), .B(new_n564), .C1(new_n568), .C2(new_n558), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n557), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G217), .B1(new_n390), .B2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT68), .ZN(new_n572));
  NAND2_X1  g386(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n194), .A2(KEYINPUT24), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT24), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G110), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n574), .B2(new_n576), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n205), .A2(G128), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n242), .A2(G119), .ZN(new_n581));
  OAI22_X1  g395(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n583), .A2(KEYINPUT23), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n242), .A2(G119), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(KEYINPUT23), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n589), .A3(new_n194), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n582), .A2(new_n590), .A3(KEYINPUT75), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT75), .B1(new_n582), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n459), .B1(new_n470), .B2(new_n237), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n194), .B1(new_n586), .B2(new_n589), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n575), .A2(G110), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n194), .A2(KEYINPUT24), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT69), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n580), .A2(new_n581), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n599), .A2(KEYINPUT70), .A3(new_n600), .A4(new_n601), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n596), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n478), .A2(KEYINPUT74), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT74), .B1(new_n478), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n595), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT77), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT74), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n604), .A2(new_n605), .ZN(new_n617));
  INV_X1    g431(.A(new_n596), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n471), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n478), .A2(new_n606), .A3(KEYINPUT74), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n595), .A3(new_n613), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n615), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n573), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(G902), .B(new_n625), .C1(new_n615), .C2(new_n623), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n572), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n613), .B1(new_n622), .B2(new_n595), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n614), .B(new_n594), .C1(new_n620), .C2(new_n621), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n572), .A2(G902), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n570), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n524), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G101), .ZN(G3));
  OAI21_X1  g454(.A(G472), .B1(new_n563), .B2(G902), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n564), .B1(new_n568), .B2(new_n558), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n629), .A2(new_n641), .A3(new_n642), .A4(new_n636), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n388), .ZN(new_n644));
  INV_X1    g458(.A(new_n396), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n310), .A2(new_n312), .ZN(new_n646));
  INV_X1    g460(.A(new_n295), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n314), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n319), .A2(new_n295), .A3(new_n316), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n323), .B(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n502), .B1(new_n521), .B2(new_n520), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n440), .A2(KEYINPUT33), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n438), .B2(new_n439), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n654), .A3(new_n435), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n435), .A2(new_n294), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n434), .B2(G478), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n644), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND2_X1  g478(.A1(new_n437), .A2(new_n441), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n665), .B(new_n502), .C1(new_n521), .C2(new_n520), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n650), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n644), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT97), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(G9));
  NOR2_X1   g485(.A1(new_n613), .A2(KEYINPUT36), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n609), .A2(KEYINPUT98), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n622), .A2(new_n674), .A3(new_n595), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n673), .A2(new_n675), .A3(new_n672), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n634), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n625), .B1(new_n632), .B2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n624), .A2(new_n626), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n573), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n679), .B1(new_n682), .B2(new_n572), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n641), .A2(new_n642), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n524), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT37), .B(G110), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n323), .B1(new_n648), .B2(new_n649), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n518), .A2(new_n519), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT20), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n518), .A2(new_n503), .A3(new_n519), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(G900), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n394), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n392), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(new_n665), .A3(new_n502), .A4(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n690), .B1(new_n691), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n666), .ZN(new_n701));
  INV_X1    g515(.A(new_n323), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n646), .A2(new_n647), .A3(new_n314), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n316), .B1(new_n319), .B2(new_n295), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n701), .A2(new_n705), .A3(KEYINPUT100), .A4(new_n698), .ZN(new_n706));
  INV_X1    g520(.A(new_n388), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n566), .A2(new_n569), .ZN(new_n708));
  INV_X1    g522(.A(new_n557), .ZN(new_n709));
  INV_X1    g523(.A(new_n679), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(new_n629), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n706), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  NAND2_X1  g527(.A1(new_n322), .A2(new_n326), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT38), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n698), .B(KEYINPUT39), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n388), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT40), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n651), .A2(new_n665), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n553), .A2(new_n544), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n532), .A2(new_n535), .A3(new_n544), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n294), .ZN(new_n723));
  OAI21_X1  g537(.A(G472), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n708), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n323), .A3(new_n683), .ZN(new_n726));
  OR4_X1    g540(.A1(new_n715), .A2(new_n719), .A3(new_n720), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G143), .ZN(G45));
  NAND3_X1  g542(.A1(new_n651), .A2(new_n659), .A3(new_n698), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n691), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n711), .A3(new_n707), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  INV_X1    g546(.A(new_n379), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n371), .B1(new_n370), .B2(new_n358), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n382), .B(new_n294), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT80), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n380), .A2(new_n382), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n387), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n661), .A2(new_n638), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  NAND3_X1  g558(.A1(new_n667), .A2(new_n638), .A3(new_n741), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT101), .B(G116), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G18));
  NOR2_X1   g561(.A1(new_n691), .A2(new_n740), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n522), .A2(new_n396), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n711), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  NAND4_X1  g565(.A1(new_n738), .A2(new_n387), .A3(new_n645), .A4(new_n739), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n643), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n691), .A2(new_n720), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT102), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT102), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  INV_X1    g574(.A(new_n729), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n748), .A2(new_n685), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  AOI21_X1  g577(.A(new_n702), .B1(new_n322), .B2(new_n326), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n382), .B1(new_n373), .B2(new_n294), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n736), .B2(new_n737), .ZN(new_n766));
  INV_X1    g580(.A(new_n387), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT103), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT103), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n385), .A2(new_n769), .A3(new_n387), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n729), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n764), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n566), .A2(new_n777), .A3(new_n569), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n709), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n635), .B1(new_n682), .B2(new_n572), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n764), .A2(new_n771), .A3(new_n773), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT105), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n764), .A2(new_n771), .A3(new_n638), .A4(new_n761), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n782), .A2(new_n785), .B1(new_n772), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n351), .ZN(G33));
  INV_X1    g602(.A(new_n699), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n764), .A2(new_n771), .A3(new_n638), .A4(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT106), .B(G134), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G36));
  AOI22_X1  g606(.A1(new_n693), .A2(new_n694), .B1(G475), .B2(new_n501), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n659), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n683), .B1(new_n642), .B2(new_n641), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(KEYINPUT44), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n382), .B1(new_n373), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n373), .ZN(new_n804));
  NAND2_X1  g618(.A1(G469), .A2(G902), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT46), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n805), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT107), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n738), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n387), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n813), .A2(KEYINPUT108), .A3(new_n717), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT108), .B1(new_n813), .B2(new_n717), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT44), .B1(new_n797), .B2(new_n798), .ZN(new_n816));
  INV_X1    g630(.A(new_n764), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n801), .A2(new_n814), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  XOR2_X1   g634(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n821));
  NAND2_X1  g635(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT47), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n812), .B(new_n387), .C1(KEYINPUT110), .C2(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n570), .A2(new_n764), .A3(new_n637), .A4(new_n761), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NOR3_X1   g641(.A1(new_n637), .A2(new_n702), .A3(new_n767), .ZN(new_n828));
  INV_X1    g642(.A(new_n794), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n738), .A2(new_n739), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT111), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n725), .B1(new_n830), .B2(new_n832), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n715), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n786), .A2(new_n772), .ZN(new_n837));
  INV_X1    g651(.A(new_n785), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT105), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n570), .A2(new_n637), .A3(new_n740), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n661), .B2(new_n667), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n757), .B1(new_n753), .B2(new_n754), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n705), .A2(new_n665), .A3(new_n651), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n844), .A2(new_n643), .A3(new_n752), .A4(KEYINPUT102), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n842), .B(new_n750), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n790), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n771), .A2(new_n685), .A3(new_n761), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  INV_X1    g663(.A(new_n698), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n522), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n793), .A2(KEYINPUT114), .A3(new_n442), .A4(new_n698), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n711), .A2(new_n851), .A3(new_n707), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n817), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n846), .A2(new_n847), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n327), .B(new_n523), .C1(new_n638), .C2(new_n685), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n327), .A2(new_n645), .A3(new_n644), .A4(new_n701), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n322), .A2(new_n323), .A3(new_n326), .A4(new_n645), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n660), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n651), .A2(new_n659), .A3(KEYINPUT112), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n859), .A2(new_n863), .A3(KEYINPUT113), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n644), .ZN(new_n866));
  INV_X1    g680(.A(new_n862), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT112), .B1(new_n651), .B2(new_n659), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n327), .A2(new_n645), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n870), .B2(KEYINPUT113), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n858), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n698), .B(KEYINPUT115), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n766), .A2(new_n767), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n754), .A2(new_n683), .A3(new_n874), .A4(new_n725), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n712), .A2(new_n731), .A3(new_n762), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n388), .A2(new_n570), .A3(new_n683), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n729), .A2(new_n683), .A3(new_n684), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n879), .A2(new_n730), .B1(new_n880), .B2(new_n748), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .A3(new_n712), .A4(new_n875), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n840), .A2(new_n855), .A3(new_n872), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n848), .A2(new_n853), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n764), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n742), .A2(new_n745), .A3(new_n750), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n759), .A4(new_n790), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n787), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n883), .A4(new_n872), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT54), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT54), .B1(new_n886), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n797), .A2(KEYINPUT116), .A3(new_n393), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n795), .A2(new_n393), .A3(new_n796), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n643), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n715), .A2(new_n702), .A3(new_n741), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(KEYINPUT50), .A3(new_n902), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n897), .A2(new_n900), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n817), .A2(new_n740), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n685), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n659), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n725), .A2(new_n637), .A3(new_n392), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n793), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n822), .A2(new_n824), .B1(new_n767), .B2(new_n832), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n901), .A2(new_n764), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n910), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n896), .B1(new_n907), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n781), .A3(new_n909), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT48), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n909), .A2(new_n912), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n389), .B1(new_n920), .B2(new_n660), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n748), .B2(new_n901), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n905), .A2(new_n906), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n914), .A2(new_n915), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n910), .A2(new_n913), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(KEYINPUT51), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n917), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n895), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n836), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT117), .B(new_n836), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G75));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n294), .B1(new_n886), .B2(new_n892), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(new_n540), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n310), .B(new_n312), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n939), .A2(new_n942), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n263), .A2(G952), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G51));
  INV_X1    g760(.A(new_n895), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n805), .B(KEYINPUT57), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n947), .A2(new_n948), .B1(new_n734), .B2(new_n733), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n938), .A2(new_n804), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G54));
  AND2_X1   g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n937), .A2(new_n518), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n518), .B1(new_n937), .B2(new_n952), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n945), .ZN(G60));
  INV_X1    g769(.A(KEYINPUT54), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT113), .B1(new_n859), .B2(new_n863), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n644), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n857), .B(new_n856), .C1(new_n958), .C2(new_n864), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n787), .A2(new_n890), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n960), .B2(new_n883), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n884), .A2(new_n885), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT54), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n656), .B(KEYINPUT59), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n652), .A2(new_n654), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n945), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n965), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT119), .B1(new_n895), .B2(new_n970), .ZN(new_n971));
  AND4_X1   g785(.A1(KEYINPUT119), .A2(new_n963), .A3(new_n964), .A4(new_n970), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT120), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n969), .B(KEYINPUT120), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G63));
  XNOR2_X1  g791(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n397), .A2(new_n294), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n886), .B2(new_n892), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n945), .B1(new_n983), .B2(new_n632), .ZN(new_n984));
  INV_X1    g798(.A(new_n678), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n985), .A2(new_n676), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n982), .A2(KEYINPUT122), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT122), .B1(new_n982), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT123), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI221_X1 g807(.A(new_n984), .B1(KEYINPUT123), .B2(KEYINPUT61), .C1(new_n988), .C2(new_n989), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G66));
  INV_X1    g809(.A(G224), .ZN(new_n996));
  OAI21_X1  g810(.A(G953), .B1(new_n395), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n959), .A2(new_n846), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n998), .B2(G953), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n318), .B(new_n300), .C1(G898), .C2(new_n263), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G69));
  NAND4_X1  g815(.A1(new_n814), .A2(new_n754), .A3(new_n815), .A4(new_n781), .ZN(new_n1002));
  AND4_X1   g816(.A1(new_n840), .A2(new_n1002), .A3(new_n790), .A4(new_n826), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n881), .A2(new_n712), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT124), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1003), .A2(new_n1005), .A3(new_n263), .A4(new_n819), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n548), .A2(new_n550), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n504), .A2(new_n506), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1007), .B(new_n1008), .Z(new_n1009));
  NAND2_X1  g823(.A1(G900), .A2(G953), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n869), .A2(new_n701), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n764), .A2(new_n638), .A3(new_n718), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n819), .A2(new_n826), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1005), .A2(new_n727), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT62), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1018));
  AOI21_X1  g832(.A(G953), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1011), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n1011), .B2(KEYINPUT125), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(G72));
  INV_X1    g839(.A(new_n721), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1017), .A2(new_n998), .A3(new_n1018), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  AOI21_X1  g843(.A(new_n1026), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n553), .A2(new_n544), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1026), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT127), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n886), .B2(new_n892), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1031), .B(KEYINPUT126), .Z(new_n1035));
  NAND4_X1  g849(.A1(new_n1003), .A2(new_n1005), .A3(new_n819), .A4(new_n998), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  NOR4_X1   g851(.A1(new_n1030), .A2(new_n945), .A3(new_n1034), .A4(new_n1037), .ZN(G57));
endmodule


