//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n205), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OR3_X1    g0016(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(G50), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n213), .A2(new_n216), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n212), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND2_X1  g0043(.A1(new_n222), .A2(G33), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  INV_X1    g0045(.A(G58), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(KEYINPUT8), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT8), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G68), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n246), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n254), .A2(G20), .B1(G150), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n251), .A2(new_n256), .B1(new_n221), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT69), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(new_n222), .A3(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n221), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(G50), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n252), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g0068(.A(new_n268), .B(KEYINPUT70), .Z(new_n269));
  NAND2_X1  g0069(.A1(new_n259), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1698), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT66), .B(G223), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n276), .B1(new_n277), .B2(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n283), .A3(G274), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(G226), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n270), .B(new_n299), .C1(G169), .C2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n259), .A2(new_n269), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n297), .A2(KEYINPUT72), .A3(G190), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n296), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n306), .A2(new_n309), .B1(G200), .B2(new_n296), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n304), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n304), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n283), .B(KEYINPUT67), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  OAI211_X1 g0117(.A(G223), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT77), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n278), .A2(KEYINPUT77), .A3(G223), .A4(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(G226), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G87), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n314), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n290), .B1(new_n232), .B2(new_n293), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n326), .A2(G179), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT78), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  INV_X1    g0130(.A(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n323), .A2(new_n324), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n320), .B2(new_n321), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n314), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT18), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n250), .A2(new_n265), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n247), .A2(new_n249), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n263), .B1(new_n261), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n273), .A2(new_n222), .A3(new_n274), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n222), .A4(new_n274), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G68), .ZN(new_n345));
  XNOR2_X1  g0145(.A(G58), .B(G68), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT16), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT76), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT7), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n340), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n316), .A2(new_n317), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n355), .B2(new_n222), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT16), .B(new_n347), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n262), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n339), .B1(new_n348), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n298), .B(new_n331), .C1(new_n333), .C2(new_n314), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n335), .A2(new_n336), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT77), .B1(new_n275), .B2(G223), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n318), .A2(new_n319), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n325), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n285), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n366), .A2(new_n329), .A3(new_n298), .A4(new_n331), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n334), .A2(new_n330), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n359), .A2(new_n361), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT18), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  INV_X1    g0172(.A(new_n339), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n357), .A2(new_n262), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n253), .B1(new_n342), .B2(new_n343), .ZN(new_n376));
  INV_X1    g0176(.A(new_n347), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n373), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(G190), .B(new_n331), .C1(new_n333), .C2(new_n314), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n334), .A2(G200), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n379), .A2(KEYINPUT79), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT79), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n327), .B1(new_n365), .B2(new_n285), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n359), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n372), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(new_n262), .A3(new_n357), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n381), .A2(new_n389), .A3(new_n339), .A4(new_n380), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(new_n372), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n371), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n253), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT68), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n244), .B(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n396), .B2(new_n277), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n262), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT11), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT11), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n400), .A3(new_n262), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n263), .A2(G68), .A3(new_n265), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n264), .A2(new_n253), .A3(G13), .A4(G20), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT12), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n399), .A2(new_n401), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT74), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n290), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G274), .ZN(new_n414));
  AND2_X1   g0214(.A1(G1), .A2(G13), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n282), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT74), .A3(new_n289), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n413), .A2(new_n417), .B1(G238), .B2(new_n294), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  OAI211_X1 g0219(.A(G226), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n420));
  OAI211_X1 g0220(.A(G232), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n420), .A2(new_n421), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n285), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n418), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n419), .B1(new_n418), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n411), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n418), .A2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n418), .A2(new_n419), .A3(new_n427), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(G179), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n411), .B1(new_n436), .B2(G169), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n410), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(G200), .B1(new_n428), .B2(new_n429), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n432), .A2(G190), .A3(new_n433), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n439), .A2(new_n440), .A3(new_n409), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT71), .ZN(new_n444));
  INV_X1    g0244(.A(G244), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n290), .B1(new_n445), .B2(new_n293), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n275), .A2(G232), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n278), .A2(G238), .A3(G1698), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n278), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n450), .B2(new_n285), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G169), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n250), .A2(new_n255), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G20), .A2(G77), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n453), .B(new_n454), .C1(new_n244), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n262), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n261), .A2(new_n277), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n263), .A2(G77), .A3(new_n265), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n444), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n451), .A2(new_n298), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n460), .B(KEYINPUT71), .C1(new_n451), .C2(G169), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n450), .A2(new_n285), .ZN(new_n466));
  INV_X1    g0266(.A(new_n446), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n468), .B2(G200), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n308), .B2(new_n468), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NOR4_X1   g0271(.A1(new_n313), .A2(new_n393), .A3(new_n443), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n288), .A2(G1), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n416), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G257), .A3(new_n283), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n479), .A2(KEYINPUT80), .A3(G257), .A4(new_n283), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT4), .A2(G244), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n315), .B(new_n485), .C1(new_n316), .C2(new_n317), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n445), .B1(new_n273), .B2(new_n274), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n486), .B(new_n487), .C1(new_n488), .C2(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g0289(.A(G250), .B1(new_n316), .B2(new_n317), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n315), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n285), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G179), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n261), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n264), .A2(G33), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n263), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n495), .A2(new_n449), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n202), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n344), .A2(G107), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n499), .B1(new_n506), .B2(new_n262), .ZN(new_n507));
  AOI21_X1  g0307(.A(G169), .B1(new_n484), .B2(new_n492), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n494), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n484), .A2(new_n308), .A3(new_n492), .ZN(new_n510));
  AOI21_X1  g0310(.A(G200), .B1(new_n484), .B2(new_n492), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT81), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n507), .B(new_n514), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n479), .A2(G270), .A3(new_n283), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n475), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G264), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n520));
  OAI211_X1 g0320(.A(G257), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n278), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n285), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n330), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n263), .A2(G116), .A3(new_n497), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n261), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n257), .A2(new_n221), .B1(G20), .B2(new_n527), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n487), .B(new_n222), .C1(G33), .C2(new_n495), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT20), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n526), .B(new_n528), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g0334(.A(KEYINPUT83), .B(KEYINPUT21), .Z(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n533), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n519), .A2(new_n524), .A3(G190), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n518), .B1(new_n285), .B2(new_n523), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n385), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n525), .A2(KEYINPUT21), .B1(new_n539), .B2(G179), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n536), .B(new_n540), .C1(new_n541), .C2(new_n537), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT82), .ZN(new_n543));
  AND3_X1   g0343(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT19), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G87), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n222), .B1(new_n547), .B2(new_n202), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n222), .B(G68), .C1(new_n316), .C2(new_n317), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n244), .B2(new_n495), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n543), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n424), .B2(new_n425), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n554), .A2(G20), .B1(G87), .B2(new_n203), .ZN(new_n555));
  INV_X1    g0355(.A(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT82), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n557), .A3(new_n262), .ZN(new_n558));
  INV_X1    g0358(.A(new_n498), .ZN(new_n559));
  INV_X1    g0359(.A(new_n455), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n455), .A2(new_n261), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G250), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n288), .B2(G1), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n264), .A2(new_n414), .A3(G45), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n283), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G238), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n285), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G179), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n330), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n563), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n285), .A2(new_n572), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n308), .A3(new_n567), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G200), .B2(new_n573), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n559), .A2(G87), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n579), .A2(new_n562), .A3(new_n558), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n542), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n516), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT85), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n222), .B(G87), .C1(new_n316), .C2(new_n317), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(KEYINPUT22), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(new_n273), .B2(new_n274), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT22), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n589), .A4(G87), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n586), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT84), .B1(new_n586), .B2(KEYINPUT22), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n587), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n222), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n449), .A2(KEYINPUT23), .A3(G20), .ZN(new_n596));
  INV_X1    g0396(.A(new_n571), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(new_n222), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n593), .A2(KEYINPUT24), .A3(new_n598), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n262), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n261), .A2(new_n449), .ZN(new_n604));
  NOR2_X1   g0404(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n604), .B2(new_n605), .ZN(new_n608));
  AOI22_X1  g0408(.A1(G107), .A2(new_n559), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n611));
  OAI211_X1 g0411(.A(G250), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n612));
  AND2_X1   g0412(.A1(KEYINPUT87), .A2(G294), .ZN(new_n613));
  NOR2_X1   g0413(.A1(KEYINPUT87), .A2(G294), .ZN(new_n614));
  OAI21_X1  g0414(.A(G33), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n285), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n474), .A2(new_n473), .B1(new_n415), .B2(new_n282), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G264), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n617), .A2(G179), .A3(new_n619), .A4(new_n475), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n285), .A2(new_n616), .B1(new_n618), .B2(G264), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n475), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT88), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT88), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n626), .A3(new_n475), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(G169), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n610), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G190), .B1(new_n625), .B2(new_n627), .ZN(new_n631));
  AOI21_X1  g0431(.A(G200), .B1(new_n623), .B2(new_n475), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n603), .B(new_n609), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n584), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n472), .A2(new_n635), .ZN(G372));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n581), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n513), .A2(new_n515), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n603), .A2(new_n609), .B1(new_n622), .B2(new_n628), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n519), .A2(new_n524), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT21), .A3(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n539), .A2(G179), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n644), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n639), .B(new_n633), .C1(new_n640), .C2(new_n646), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n494), .A2(new_n507), .A3(new_n508), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n638), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n573), .A2(new_n330), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n298), .B(new_n568), .C1(new_n285), .C2(new_n572), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT90), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n574), .B(new_n653), .C1(new_n330), .C2(new_n573), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n563), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n648), .A2(new_n582), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n637), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n472), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT91), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n468), .A2(new_n330), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT71), .B1(new_n661), .B2(new_n460), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n464), .A2(new_n463), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT92), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT92), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n462), .A2(new_n464), .A3(new_n665), .A4(new_n463), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n442), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n438), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n382), .A2(new_n387), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n391), .B1(new_n669), .B2(KEYINPUT17), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n671), .A2(new_n371), .B1(new_n312), .B2(new_n311), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n672), .A2(new_n300), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n660), .A2(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n264), .A2(new_n222), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G343), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n645), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT94), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n680), .B1(new_n603), .B2(new_n609), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n634), .A2(new_n684), .B1(new_n630), .B2(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n630), .B2(new_n681), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n537), .A2(new_n680), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT93), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n645), .A3(new_n540), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n645), .B2(new_n690), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n685), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n695), .ZN(G399));
  NOR3_X1   g0496(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n214), .A2(new_n287), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(G1), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n219), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n702), .B(new_n680), .C1(new_n649), .C2(new_n657), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n639), .A2(new_n648), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT95), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n630), .A2(new_n645), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n516), .A2(KEYINPUT95), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n655), .A2(new_n581), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(new_n633), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n656), .A2(new_n637), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n509), .A2(new_n581), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT26), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n712), .A2(new_n655), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n681), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n703), .B1(new_n716), .B2(new_n702), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n539), .A2(new_n484), .A3(new_n623), .A4(new_n492), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n574), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n484), .A2(new_n492), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n623), .A2(new_n524), .A3(new_n519), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT30), .A4(new_n651), .ZN(new_n724));
  AOI21_X1  g0524(.A(G179), .B1(new_n519), .B2(new_n524), .ZN(new_n725));
  INV_X1    g0525(.A(new_n573), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n493), .A2(new_n725), .A3(new_n624), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n721), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n681), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n630), .A2(new_n633), .A3(new_n680), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n731), .B(new_n732), .C1(new_n584), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n718), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n701), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n260), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n264), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n698), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n693), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n692), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n278), .A2(new_n214), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n214), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n239), .A2(G45), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n355), .A2(new_n214), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n220), .B2(new_n288), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n221), .B1(G20), .B2(new_n330), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n743), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n222), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n308), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n449), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n298), .A2(new_n385), .A3(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n495), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n762), .B(new_n766), .C1(G87), .C2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n222), .A2(new_n298), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(new_n385), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n278), .B1(new_n771), .B2(new_n246), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(G77), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n760), .A2(new_n773), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n770), .A2(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n308), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(G190), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G50), .A2(new_n782), .B1(new_n783), .B2(G68), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n769), .A2(new_n776), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n767), .B(KEYINPUT96), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n522), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n613), .A2(new_n614), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n765), .A2(new_n789), .B1(new_n761), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G326), .B2(new_n782), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(new_n783), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n278), .B1(new_n775), .B2(G311), .ZN(new_n798));
  INV_X1    g0598(.A(new_n771), .ZN(new_n799));
  INV_X1    g0599(.A(new_n777), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G322), .B1(new_n800), .B2(G329), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n785), .B1(new_n788), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT98), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n756), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n759), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n755), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n692), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n745), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n658), .A2(new_n680), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n460), .A2(new_n681), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n664), .A2(new_n666), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n465), .A2(new_n470), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n813), .B(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n743), .B1(new_n820), .B2(new_n735), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n735), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n756), .A2(new_n753), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n743), .B1(G77), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n799), .A2(G143), .B1(new_n775), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(new_n782), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  INV_X1    g0629(.A(new_n783), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n826), .B1(new_n827), .B2(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n786), .A2(G50), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n278), .B1(new_n777), .B2(new_n836), .C1(new_n253), .C2(new_n761), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G58), .B2(new_n764), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n827), .A2(new_n522), .B1(new_n774), .B2(new_n527), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n840), .B1(new_n844), .B2(G283), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT100), .Z(new_n846));
  AOI211_X1 g0646(.A(new_n278), .B(new_n766), .C1(G294), .C2(new_n799), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n761), .A2(new_n547), .B1(new_n777), .B2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT101), .Z(new_n850));
  OAI211_X1 g0650(.A(new_n847), .B(new_n850), .C1(new_n449), .C2(new_n787), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n839), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n825), .B1(new_n852), .B2(new_n756), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n754), .B2(new_n818), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n822), .A2(new_n854), .ZN(G384));
  XOR2_X1   g0655(.A(new_n503), .B(KEYINPUT102), .Z(new_n856));
  INV_X1    g0656(.A(KEYINPUT35), .ZN(new_n857));
  OAI211_X1 g0657(.A(G116), .B(new_n223), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n277), .B(new_n219), .C1(G58), .C2(G68), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n252), .B2(G68), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n264), .B(G13), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n410), .A2(new_n681), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n438), .A2(new_n442), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(G169), .B1(new_n428), .B2(new_n429), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT14), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n434), .A3(new_n430), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n410), .B(new_n681), .C1(new_n871), .C2(new_n441), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n868), .A2(new_n872), .B1(new_n816), .B2(new_n817), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n732), .B1(new_n584), .B2(new_n733), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT105), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n728), .A2(new_n875), .A3(new_n681), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n728), .B2(new_n681), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT31), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n873), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT106), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n340), .A2(KEYINPUT7), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(G68), .C1(new_n340), .C2(new_n353), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT16), .B1(new_n884), .B2(new_n347), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n339), .B1(new_n358), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n679), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n362), .A2(new_n370), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n670), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n886), .A2(new_n361), .A3(new_n367), .A4(new_n368), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n382), .A2(new_n387), .A3(new_n890), .A4(new_n887), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n382), .A2(new_n387), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT37), .B1(new_n359), .B2(new_n679), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n369), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(KEYINPUT37), .A2(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n882), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n382), .A2(new_n387), .A3(new_n369), .A4(new_n893), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT38), .B(new_n899), .C1(new_n392), .C2(new_n887), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n873), .B(KEYINPUT106), .C1(new_n874), .C2(new_n878), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n881), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n359), .A2(new_n679), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n670), .B2(new_n888), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n369), .A2(new_n390), .A3(new_n906), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n892), .A2(new_n894), .B1(KEYINPUT37), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n882), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n900), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n873), .B(KEYINPUT40), .C1(new_n874), .C2(new_n878), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n905), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n472), .B1(new_n874), .B2(new_n878), .ZN(new_n914));
  OAI21_X1  g0714(.A(G330), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n871), .A2(new_n410), .A3(new_n680), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n919));
  AND3_X1   g0719(.A1(new_n910), .A2(new_n900), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n896), .B2(new_n900), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n868), .A2(new_n872), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n680), .B(new_n818), .C1(new_n649), .C2(new_n657), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n465), .A2(new_n681), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n901), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n888), .A2(new_n679), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n923), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n717), .A2(new_n472), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n673), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n916), .A2(new_n936), .B1(new_n264), .B2(new_n739), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n916), .A2(new_n936), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n866), .B1(new_n937), .B2(new_n938), .ZN(G367));
  NAND3_X1  g0739(.A1(new_n558), .A2(new_n562), .A3(new_n580), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n681), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n709), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n655), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n706), .B(new_n708), .C1(new_n507), .C2(new_n680), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n509), .A2(new_n681), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT42), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(new_n950), .A3(new_n685), .A4(new_n683), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT108), .ZN(new_n952));
  INV_X1    g0752(.A(new_n949), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT42), .B1(new_n953), .B2(new_n686), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n509), .B1(new_n949), .B2(new_n640), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n954), .B1(new_n681), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n945), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n694), .A2(new_n949), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT109), .Z(new_n959));
  OR2_X1    g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n959), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT43), .B2(new_n944), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n698), .B(KEYINPUT41), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT110), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n688), .A2(new_n967), .A3(new_n949), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT110), .B1(new_n953), .B2(new_n687), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n953), .A2(new_n687), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT45), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n695), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n686), .A2(KEYINPUT112), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(new_n693), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n683), .A2(new_n685), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n737), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n977), .A2(new_n978), .A3(new_n694), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n980), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n966), .B1(new_n990), .B2(new_n737), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n963), .B(new_n965), .C1(new_n991), .C2(new_n741), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n230), .A2(new_n214), .A3(new_n355), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n757), .B1(new_n214), .B2(new_n455), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n743), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n844), .A2(G159), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n774), .A2(new_n252), .B1(new_n777), .B2(new_n828), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n355), .B(new_n997), .C1(G150), .C2(new_n799), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n761), .A2(new_n277), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G68), .B2(new_n764), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n782), .A2(G143), .B1(new_n768), .B2(G58), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n827), .A2(new_n848), .B1(new_n761), .B2(new_n495), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G107), .B2(new_n764), .ZN(new_n1004));
  INV_X1    g0804(.A(G317), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n771), .A2(new_n522), .B1(new_n777), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n278), .B(new_n1006), .C1(G283), .C2(new_n775), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n767), .A2(new_n527), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1004), .B(new_n1007), .C1(KEYINPUT46), .C2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n786), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n843), .B2(new_n789), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1002), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n995), .B1(new_n1013), .B2(new_n756), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n942), .A2(new_n755), .A3(new_n943), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n992), .A2(new_n1016), .ZN(G387));
  OR2_X1    g0817(.A1(new_n685), .A2(new_n809), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n747), .A2(new_n697), .B1(G107), .B2(new_n214), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n697), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n1020), .C1(G68), .C2(G77), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n250), .A2(new_n252), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT50), .Z(new_n1023));
  AOI21_X1  g0823(.A(new_n750), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n235), .A2(G45), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1019), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n743), .B1(new_n1026), .B2(new_n758), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n771), .A2(new_n252), .B1(new_n774), .B2(new_n253), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n355), .B(new_n1028), .C1(G150), .C2(new_n800), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n783), .A2(new_n250), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n765), .A2(new_n455), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G159), .B2(new_n782), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n761), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n768), .A2(G77), .B1(new_n1033), .B2(G97), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n278), .B1(new_n800), .B2(G326), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n765), .A2(new_n790), .B1(new_n789), .B2(new_n767), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT113), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n771), .A2(new_n1005), .B1(new_n774), .B2(new_n522), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G322), .B2(new_n782), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n843), .B2(new_n848), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1036), .B1(new_n527), .B2(new_n761), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1035), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT114), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n806), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1027), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n986), .A2(new_n741), .B1(new_n1018), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n987), .A2(new_n742), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n986), .A2(new_n737), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(G393));
  NAND2_X1  g0856(.A1(new_n977), .A2(new_n694), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n972), .A2(new_n975), .A3(new_n695), .A4(new_n976), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n741), .A3(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n757), .B1(new_n495), .B2(new_n214), .C1(new_n242), .C2(new_n750), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n743), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n767), .A2(new_n790), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n762), .B(new_n1062), .C1(G116), .C2(new_n764), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n800), .A2(G322), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n278), .B(new_n1064), .C1(G294), .C2(new_n775), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(new_n843), .C2(new_n522), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G317), .A2(new_n782), .B1(new_n799), .B2(G311), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G150), .A2(new_n782), .B1(new_n799), .B2(G159), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1069), .B(new_n1070), .Z(new_n1071));
  INV_X1    g0871(.A(G143), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n278), .B1(new_n777), .B2(new_n1072), .C1(new_n338), .C2(new_n774), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n765), .A2(new_n277), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n253), .A2(new_n767), .B1(new_n761), .B2(new_n547), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n843), .B2(new_n252), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1066), .A2(new_n1068), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1061), .B1(new_n1078), .B2(new_n756), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n949), .B2(new_n809), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1059), .A2(KEYINPUT116), .A3(new_n1080), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n698), .B1(new_n1085), .B2(new_n987), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1083), .A2(new_n1084), .B1(new_n990), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  NOR2_X1   g0888(.A1(new_n516), .A2(KEYINPUT95), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n705), .B(new_n509), .C1(new_n513), .C2(new_n515), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n709), .B(new_n633), .C1(new_n640), .C2(new_n646), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n712), .A2(new_n655), .A3(new_n714), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n680), .B(new_n818), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n734), .A2(G330), .A3(new_n818), .A4(new_n924), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1094), .A2(new_n928), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(G330), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n874), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n878), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n818), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n925), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n925), .B1(new_n735), .B2(new_n819), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n873), .B(G330), .C1(new_n874), .C2(new_n878), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n926), .A2(new_n928), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1096), .A2(new_n1102), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n472), .A2(new_n1100), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n934), .A2(new_n673), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n922), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n910), .A2(new_n900), .A3(new_n919), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(new_n929), .C2(new_n918), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n918), .B1(new_n910), .B2(new_n900), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n927), .B1(new_n716), .B2(new_n818), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n925), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1114), .A2(new_n1117), .A3(new_n1095), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1104), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1111), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1104), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1114), .A2(new_n1117), .A3(new_n1095), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1110), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n742), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1112), .A2(new_n753), .A3(new_n1113), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n743), .B1(new_n250), .B2(new_n824), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT117), .Z(new_n1130));
  AOI21_X1  g0930(.A(new_n355), .B1(new_n800), .B2(G125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n836), .B2(new_n771), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT53), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n767), .A2(new_n829), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT118), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1135), .B1(new_n1133), .B2(new_n1134), .C1(new_n774), .C2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1033), .A2(G50), .B1(new_n764), .B2(G159), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n827), .C1(new_n843), .C2(new_n828), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1074), .B1(G68), .B2(new_n1033), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n278), .B1(new_n775), .B2(G97), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n799), .A2(G116), .B1(new_n800), .B2(G294), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n782), .A2(G283), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n843), .A2(new_n449), .B1(new_n547), .B2(new_n787), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1139), .A2(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n1149), .B2(new_n756), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT119), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1127), .A2(new_n741), .B1(new_n1128), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1126), .A2(new_n1152), .ZN(G378));
  AOI21_X1  g0953(.A(new_n1109), .B1(new_n1127), .B2(new_n1110), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n923), .A2(new_n930), .A3(new_n932), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n879), .A2(new_n880), .B1(new_n896), .B2(new_n900), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT40), .B1(new_n1156), .B2(new_n902), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n270), .A2(new_n679), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n313), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n300), .B(new_n1158), .C1(new_n311), .C2(new_n312), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(G330), .B1(new_n911), .B2(new_n912), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1157), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1163), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n912), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n910), .A2(new_n900), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1097), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1172), .B1(new_n905), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1155), .B1(new_n1169), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1167), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n905), .A2(new_n1175), .A3(new_n1172), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n933), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1109), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1125), .A2(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n933), .A2(new_n1179), .A3(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n931), .B1(new_n1186), .B2(new_n918), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1178), .A2(new_n1179), .B1(new_n1187), .B2(new_n930), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT124), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1184), .A2(new_n1189), .A3(new_n1190), .A4(KEYINPUT57), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n698), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT122), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1155), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT123), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1178), .A2(new_n1179), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT123), .B1(new_n1169), .B2(new_n1176), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1194), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1178), .A2(new_n1179), .A3(new_n1195), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1198), .A2(new_n1202), .B1(new_n1183), .B2(new_n1125), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT125), .B1(new_n1203), .B2(KEYINPUT57), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1196), .A2(new_n1197), .A3(new_n1194), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1200), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1184), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT125), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1192), .A2(new_n1204), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n743), .B1(G50), .B2(new_n824), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT121), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1167), .A2(new_n754), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(G33), .A2(G41), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G50), .B(new_n1215), .C1(new_n355), .C2(new_n287), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n830), .A2(new_n495), .B1(new_n246), .B2(new_n761), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G116), .B2(new_n782), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G41), .B(new_n278), .C1(new_n800), .C2(G283), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n799), .A2(G107), .B1(new_n775), .B2(new_n560), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n768), .A2(G77), .B1(new_n764), .B2(G68), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n771), .A2(new_n1141), .B1(new_n774), .B2(new_n828), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G150), .B2(new_n764), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G125), .A2(new_n782), .B1(new_n783), .B2(G132), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n1138), .C2(new_n767), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1230));
  INV_X1    g1030(.A(G124), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1215), .B1(new_n777), .B2(new_n1231), .C1(new_n778), .C2(new_n761), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT120), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1224), .B1(new_n1223), .B2(new_n1222), .C1(new_n1229), .C2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1213), .B(new_n1214), .C1(new_n756), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n741), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1211), .A2(new_n1238), .ZN(G375));
  INV_X1    g1039(.A(new_n1107), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n925), .A2(new_n753), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n743), .B1(G68), .B2(new_n824), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n844), .A2(new_n1137), .B1(G159), .B2(new_n786), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n771), .A2(new_n828), .B1(new_n777), .B2(new_n1141), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n355), .B(new_n1244), .C1(G150), .C2(new_n775), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n827), .A2(new_n836), .B1(new_n761), .B2(new_n246), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G50), .B2(new_n764), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n844), .A2(G116), .B1(G97), .B2(new_n786), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n771), .A2(new_n790), .B1(new_n777), .B2(new_n522), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n278), .B(new_n1250), .C1(G107), .C2(new_n775), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n999), .B(new_n1031), .C1(G294), .C2(new_n782), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1242), .B1(new_n1254), .B2(new_n756), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1240), .A2(new_n741), .B1(new_n1241), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1110), .A2(new_n966), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1240), .A2(new_n1183), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1258), .B2(new_n1259), .ZN(G381));
  NAND3_X1  g1060(.A1(new_n992), .A2(new_n1016), .A3(new_n1087), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n811), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1262));
  OR3_X1    g1062(.A1(new_n1262), .A2(KEYINPUT126), .A3(G384), .ZN(new_n1263));
  INV_X1    g1063(.A(G381), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT126), .B1(new_n1262), .B2(G384), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G378), .A2(new_n1261), .A3(G375), .A4(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  INV_X1    g1068(.A(G343), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1211), .A2(G378), .A3(new_n1238), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1236), .B1(new_n1189), .B2(new_n741), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1207), .B2(new_n966), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1268), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1271), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1259), .A2(new_n1280), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1240), .A2(new_n1183), .A3(KEYINPUT60), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n742), .B(new_n1111), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(G384), .A3(new_n1256), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1283), .B2(new_n1256), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1271), .A2(G2897), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G2897), .B(new_n1271), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1274), .B1(new_n1279), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1270), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1287), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n965), .A2(new_n963), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n990), .A2(new_n737), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n966), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1302), .B2(new_n740), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1016), .ZN(new_n1304));
  OAI21_X1  g1104(.A(G390), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1306), .A2(KEYINPUT127), .A3(new_n1262), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1262), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1305), .B(new_n1261), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1261), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1087), .B1(new_n992), .B2(new_n1016), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1309), .B1(new_n1312), .B2(new_n1307), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1279), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1293), .A2(new_n1298), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1279), .A2(new_n1316), .A3(new_n1287), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1279), .B2(new_n1287), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1317), .A2(new_n1292), .A3(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1315), .B1(new_n1319), .B2(new_n1313), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1268), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1275), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1287), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1297), .A3(new_n1275), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1325), .A2(new_n1313), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1313), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


