

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723;

  NAND2_X1 U368 ( .A1(n399), .A2(n420), .ZN(n347) );
  OR2_X1 U369 ( .A1(n672), .A2(n409), .ZN(n408) );
  XNOR2_X1 U370 ( .A(n562), .B(n402), .ZN(n590) );
  OR2_X1 U371 ( .A1(n608), .A2(G902), .ZN(n417) );
  INV_X1 U372 ( .A(G143), .ZN(n413) );
  INV_X1 U373 ( .A(KEYINPUT3), .ZN(n458) );
  XNOR2_X2 U374 ( .A(n346), .B(KEYINPUT71), .ZN(n586) );
  NAND2_X2 U375 ( .A1(n395), .A2(n567), .ZN(n346) );
  XNOR2_X2 U376 ( .A(n347), .B(n419), .ZN(n718) );
  XNOR2_X2 U377 ( .A(n348), .B(n376), .ZN(n696) );
  XNOR2_X2 U378 ( .A(n473), .B(n501), .ZN(n348) );
  XNOR2_X2 U379 ( .A(n514), .B(n433), .ZN(n708) );
  XNOR2_X2 U380 ( .A(n475), .B(n412), .ZN(n514) );
  BUF_X2 U381 ( .A(n687), .Z(n691) );
  INV_X1 U382 ( .A(n590), .ZN(n651) );
  INV_X1 U383 ( .A(G953), .ZN(n710) );
  NOR2_X2 U384 ( .A1(n349), .A2(n598), .ZN(n599) );
  XNOR2_X2 U385 ( .A(n361), .B(n537), .ZN(n719) );
  XNOR2_X2 U386 ( .A(n403), .B(n456), .ZN(n562) );
  INV_X1 U387 ( .A(KEYINPUT16), .ZN(n377) );
  NOR2_X1 U388 ( .A1(n655), .A2(n540), .ZN(n610) );
  INV_X1 U389 ( .A(n635), .ZN(n597) );
  NOR2_X2 U390 ( .A1(G902), .A2(n685), .ZN(n509) );
  XNOR2_X1 U391 ( .A(n474), .B(n377), .ZN(n376) );
  XNOR2_X1 U392 ( .A(n378), .B(G110), .ZN(n474) );
  XNOR2_X1 U393 ( .A(n483), .B(n397), .ZN(n707) );
  XNOR2_X1 U394 ( .A(n368), .B(n541), .ZN(n349) );
  XNOR2_X1 U395 ( .A(n368), .B(n541), .ZN(n702) );
  XOR2_X1 U396 ( .A(G146), .B(G125), .Z(n483) );
  INV_X1 U397 ( .A(G137), .ZN(n431) );
  XNOR2_X1 U398 ( .A(G131), .B(KEYINPUT4), .ZN(n432) );
  OR2_X1 U399 ( .A1(n455), .A2(G902), .ZN(n403) );
  INV_X1 U400 ( .A(KEYINPUT19), .ZN(n491) );
  NOR2_X1 U401 ( .A1(n610), .A2(n350), .ZN(n389) );
  XNOR2_X1 U402 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U403 ( .A(n708), .B(G146), .ZN(n461) );
  INV_X1 U404 ( .A(KEYINPUT1), .ZN(n402) );
  XOR2_X1 U405 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n497) );
  NOR2_X1 U406 ( .A1(G953), .A2(G237), .ZN(n498) );
  XNOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT8), .ZN(n448) );
  XNOR2_X1 U408 ( .A(KEYINPUT69), .B(KEYINPUT38), .ZN(n411) );
  XOR2_X1 U409 ( .A(n454), .B(n453), .Z(n533) );
  NAND2_X1 U410 ( .A1(n460), .A2(n459), .ZN(n381) );
  INV_X1 U411 ( .A(G119), .ZN(n378) );
  XNOR2_X1 U412 ( .A(G137), .B(G128), .ZN(n445) );
  XNOR2_X1 U413 ( .A(KEYINPUT10), .B(G140), .ZN(n397) );
  NAND2_X1 U414 ( .A1(n625), .A2(n551), .ZN(n592) );
  NOR2_X1 U415 ( .A1(n559), .A2(n550), .ZN(n551) );
  NOR2_X1 U416 ( .A1(n559), .A2(n384), .ZN(n561) );
  XOR2_X1 U417 ( .A(G475), .B(n510), .Z(n528) );
  XNOR2_X1 U418 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U419 ( .A(KEYINPUT83), .ZN(n422) );
  NAND2_X1 U420 ( .A1(n550), .A2(n590), .ZN(n407) );
  XNOR2_X1 U421 ( .A(n461), .B(n434), .ZN(n455) );
  INV_X1 U422 ( .A(KEYINPUT40), .ZN(n414) );
  NAND2_X1 U423 ( .A1(n596), .A2(n625), .ZN(n415) );
  XNOR2_X1 U424 ( .A(n720), .B(KEYINPUT78), .ZN(n392) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n390) );
  XOR2_X1 U426 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n503) );
  XNOR2_X1 U427 ( .A(G143), .B(KEYINPUT95), .ZN(n502) );
  XNOR2_X1 U428 ( .A(G113), .B(G131), .ZN(n496) );
  XNOR2_X1 U429 ( .A(n709), .B(KEYINPUT70), .ZN(n598) );
  XOR2_X1 U430 ( .A(G107), .B(KEYINPUT67), .Z(n482) );
  XNOR2_X1 U431 ( .A(KEYINPUT84), .B(KEYINPUT18), .ZN(n478) );
  NAND2_X1 U432 ( .A1(G234), .A2(G237), .ZN(n466) );
  XNOR2_X1 U433 ( .A(G902), .B(KEYINPUT15), .ZN(n600) );
  OR2_X1 U434 ( .A1(G237), .A2(G902), .ZN(n487) );
  INV_X1 U435 ( .A(KEYINPUT30), .ZN(n570) );
  NOR2_X1 U436 ( .A1(n654), .A2(n533), .ZN(n650) );
  XNOR2_X1 U437 ( .A(G116), .B(G107), .ZN(n511) );
  INV_X1 U438 ( .A(G134), .ZN(n412) );
  XNOR2_X1 U439 ( .A(G101), .B(G104), .ZN(n425) );
  XOR2_X1 U440 ( .A(G140), .B(G110), .Z(n426) );
  XNOR2_X1 U441 ( .A(n588), .B(n587), .ZN(n596) );
  AND2_X1 U442 ( .A1(n572), .A2(n568), .ZN(n395) );
  XNOR2_X1 U443 ( .A(n571), .B(n570), .ZN(n572) );
  INV_X1 U444 ( .A(n409), .ZN(n585) );
  AND2_X1 U445 ( .A1(n650), .A2(n562), .ZN(n567) );
  XNOR2_X1 U446 ( .A(n461), .B(n418), .ZN(n608) );
  XNOR2_X1 U447 ( .A(n464), .B(n473), .ZN(n418) );
  XNOR2_X1 U448 ( .A(n452), .B(n396), .ZN(n693) );
  XNOR2_X1 U449 ( .A(n707), .B(n447), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n636), .B(n369), .ZN(n678) );
  XNOR2_X1 U451 ( .A(n370), .B(KEYINPUT2), .ZN(n369) );
  INV_X1 U452 ( .A(KEYINPUT76), .ZN(n370) );
  INV_X1 U453 ( .A(KEYINPUT42), .ZN(n416) );
  INV_X1 U454 ( .A(KEYINPUT35), .ZN(n419) );
  INV_X1 U455 ( .A(n574), .ZN(n420) );
  INV_X1 U456 ( .A(n662), .ZN(n383) );
  AND2_X1 U457 ( .A1(n528), .A2(n524), .ZN(n522) );
  XNOR2_X1 U458 ( .A(n406), .B(n405), .ZN(n540) );
  INV_X1 U459 ( .A(KEYINPUT80), .ZN(n405) );
  INV_X1 U460 ( .A(KEYINPUT60), .ZN(n363) );
  XNOR2_X1 U461 ( .A(n605), .B(n357), .ZN(n606) );
  INV_X1 U462 ( .A(KEYINPUT56), .ZN(n365) );
  AND2_X1 U463 ( .A1(n523), .A2(n558), .ZN(n350) );
  XOR2_X1 U464 ( .A(KEYINPUT68), .B(n465), .Z(n351) );
  XOR2_X1 U465 ( .A(n483), .B(n482), .Z(n352) );
  NOR2_X1 U466 ( .A1(n641), .A2(n654), .ZN(n353) );
  AND2_X1 U467 ( .A1(n718), .A2(n618), .ZN(n354) );
  AND2_X1 U468 ( .A1(n597), .A2(n634), .ZN(n355) );
  XOR2_X1 U469 ( .A(n422), .B(KEYINPUT0), .Z(n356) );
  XNOR2_X1 U470 ( .A(n455), .B(n437), .ZN(n357) );
  XOR2_X1 U471 ( .A(n685), .B(n684), .Z(n358) );
  XOR2_X1 U472 ( .A(n608), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U473 ( .A(n682), .B(n424), .Z(n360) );
  NOR2_X1 U474 ( .A1(G952), .A2(n710), .ZN(n695) );
  INV_X1 U475 ( .A(n695), .ZN(n373) );
  NOR2_X2 U476 ( .A1(n539), .A2(n536), .ZN(n361) );
  XNOR2_X1 U477 ( .A(n362), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U478 ( .A1(n372), .A2(n373), .ZN(n362) );
  XNOR2_X1 U479 ( .A(n364), .B(n363), .ZN(G60) );
  NAND2_X1 U480 ( .A1(n371), .A2(n373), .ZN(n364) );
  XNOR2_X1 U481 ( .A(n366), .B(n365), .ZN(G51) );
  NAND2_X1 U482 ( .A1(n374), .A2(n373), .ZN(n366) );
  XNOR2_X1 U483 ( .A(n707), .B(n500), .ZN(n507) );
  XNOR2_X1 U484 ( .A(n507), .B(n506), .ZN(n685) );
  NAND2_X1 U485 ( .A1(n388), .A2(n354), .ZN(n387) );
  INV_X2 U486 ( .A(n569), .ZN(n384) );
  NAND2_X1 U487 ( .A1(n563), .A2(n562), .ZN(n409) );
  XNOR2_X1 U488 ( .A(n387), .B(n538), .ZN(n386) );
  NAND2_X1 U489 ( .A1(n564), .A2(n492), .ZN(n493) );
  XNOR2_X1 U490 ( .A(n552), .B(n491), .ZN(n564) );
  NAND2_X1 U491 ( .A1(n386), .A2(n389), .ZN(n368) );
  XNOR2_X1 U492 ( .A(n686), .B(n358), .ZN(n371) );
  XNOR2_X1 U493 ( .A(n609), .B(n359), .ZN(n372) );
  XNOR2_X1 U494 ( .A(n683), .B(n360), .ZN(n374) );
  XNOR2_X1 U495 ( .A(n375), .B(KEYINPUT46), .ZN(n394) );
  NOR2_X2 U496 ( .A1(n722), .A2(n723), .ZN(n375) );
  XNOR2_X1 U497 ( .A(n499), .B(n423), .ZN(n500) );
  INV_X1 U498 ( .A(n673), .ZN(n382) );
  XNOR2_X2 U499 ( .A(n381), .B(n380), .ZN(n473) );
  XNOR2_X2 U500 ( .A(G116), .B(G113), .ZN(n380) );
  AND2_X2 U501 ( .A1(n385), .A2(n353), .ZN(n421) );
  NAND2_X1 U502 ( .A1(n385), .A2(n382), .ZN(n401) );
  AND2_X1 U503 ( .A1(n385), .A2(n383), .ZN(n495) );
  AND2_X1 U504 ( .A1(n385), .A2(n384), .ZN(n494) );
  XNOR2_X2 U505 ( .A(n493), .B(n356), .ZN(n385) );
  INV_X1 U506 ( .A(n719), .ZN(n388) );
  XNOR2_X2 U507 ( .A(n391), .B(n390), .ZN(n410) );
  NAND2_X1 U508 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X2 U509 ( .A(n557), .B(KEYINPUT108), .ZN(n720) );
  AND2_X1 U510 ( .A1(n394), .A2(n589), .ZN(n393) );
  NAND2_X1 U511 ( .A1(n586), .A2(n638), .ZN(n588) );
  XNOR2_X1 U512 ( .A(n401), .B(n400), .ZN(n399) );
  INV_X1 U513 ( .A(KEYINPUT34), .ZN(n400) );
  NOR2_X1 U514 ( .A1(n702), .A2(n709), .ZN(n636) );
  XNOR2_X2 U515 ( .A(n404), .B(n490), .ZN(n552) );
  NAND2_X1 U516 ( .A1(n595), .A2(n637), .ZN(n404) );
  XNOR2_X2 U517 ( .A(n489), .B(n488), .ZN(n595) );
  NOR2_X1 U518 ( .A1(n539), .A2(n407), .ZN(n406) );
  XNOR2_X2 U519 ( .A(n421), .B(n530), .ZN(n539) );
  NAND2_X2 U520 ( .A1(n410), .A2(n355), .ZN(n709) );
  XNOR2_X2 U521 ( .A(n408), .B(n416), .ZN(n723) );
  XNOR2_X1 U522 ( .A(n584), .B(KEYINPUT41), .ZN(n672) );
  XNOR2_X1 U523 ( .A(n595), .B(n411), .ZN(n638) );
  XNOR2_X2 U524 ( .A(n413), .B(G128), .ZN(n475) );
  INV_X1 U525 ( .A(n672), .ZN(n666) );
  XNOR2_X2 U526 ( .A(n415), .B(n414), .ZN(n722) );
  XNOR2_X2 U527 ( .A(n417), .B(n351), .ZN(n569) );
  NAND2_X1 U528 ( .A1(n606), .A2(n373), .ZN(n607) );
  XOR2_X2 U529 ( .A(n384), .B(KEYINPUT6), .Z(n550) );
  AND2_X1 U530 ( .A1(G214), .A2(n498), .ZN(n423) );
  XNOR2_X1 U531 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n424) );
  INV_X1 U532 ( .A(KEYINPUT44), .ZN(n538) );
  XNOR2_X1 U533 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U534 ( .A(n484), .B(n352), .ZN(n485) );
  INV_X1 U535 ( .A(KEYINPUT82), .ZN(n490) );
  XNOR2_X1 U536 ( .A(n486), .B(n485), .ZN(n682) );
  XNOR2_X1 U537 ( .A(KEYINPUT36), .B(KEYINPUT81), .ZN(n554) );
  INV_X1 U538 ( .A(KEYINPUT59), .ZN(n684) );
  XNOR2_X1 U539 ( .A(n555), .B(n554), .ZN(n556) );
  INV_X1 U540 ( .A(n482), .ZN(n428) );
  XNOR2_X1 U541 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U542 ( .A(n428), .B(n427), .ZN(n430) );
  NAND2_X1 U543 ( .A1(G227), .A2(n710), .ZN(n429) );
  XNOR2_X1 U544 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U545 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n436) );
  XNOR2_X1 U546 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n435) );
  XNOR2_X1 U547 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U548 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n440) );
  NAND2_X1 U549 ( .A1(G234), .A2(n600), .ZN(n438) );
  XNOR2_X1 U550 ( .A(KEYINPUT20), .B(n438), .ZN(n441) );
  NAND2_X1 U551 ( .A1(G221), .A2(n441), .ZN(n439) );
  XNOR2_X1 U552 ( .A(n440), .B(n439), .ZN(n654) );
  XOR2_X1 U553 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n443) );
  NAND2_X1 U554 ( .A1(G217), .A2(n441), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U556 ( .A(KEYINPUT25), .B(n444), .ZN(n454) );
  XOR2_X1 U557 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n446) );
  XNOR2_X1 U558 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U559 ( .A(n474), .B(KEYINPUT23), .Z(n451) );
  NAND2_X1 U560 ( .A1(n710), .A2(G234), .ZN(n449) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n515) );
  NAND2_X1 U562 ( .A1(G221), .A2(n515), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n450), .B(n451), .ZN(n452) );
  NOR2_X1 U564 ( .A1(G902), .A2(n693), .ZN(n453) );
  XNOR2_X1 U565 ( .A(KEYINPUT66), .B(G469), .ZN(n456) );
  INV_X1 U566 ( .A(G101), .ZN(n457) );
  NAND2_X1 U567 ( .A1(n457), .A2(KEYINPUT3), .ZN(n460) );
  NAND2_X1 U568 ( .A1(n458), .A2(G101), .ZN(n459) );
  XOR2_X1 U569 ( .A(G119), .B(KEYINPUT5), .Z(n463) );
  NAND2_X1 U570 ( .A1(n498), .A2(G210), .ZN(n462) );
  XOR2_X1 U571 ( .A(n463), .B(n462), .Z(n464) );
  XOR2_X1 U572 ( .A(G472), .B(KEYINPUT94), .Z(n465) );
  XNOR2_X1 U573 ( .A(n466), .B(KEYINPUT14), .ZN(n468) );
  NAND2_X1 U574 ( .A1(n468), .A2(G952), .ZN(n467) );
  XNOR2_X1 U575 ( .A(n467), .B(KEYINPUT86), .ZN(n671) );
  NOR2_X1 U576 ( .A1(G953), .A2(n671), .ZN(n545) );
  NAND2_X1 U577 ( .A1(n468), .A2(G902), .ZN(n469) );
  XNOR2_X1 U578 ( .A(KEYINPUT88), .B(n469), .ZN(n542) );
  NOR2_X1 U579 ( .A1(G898), .A2(n710), .ZN(n470) );
  XNOR2_X1 U580 ( .A(KEYINPUT87), .B(n470), .ZN(n698) );
  NOR2_X1 U581 ( .A1(n542), .A2(n698), .ZN(n471) );
  NOR2_X1 U582 ( .A1(n545), .A2(n471), .ZN(n472) );
  XNOR2_X1 U583 ( .A(KEYINPUT89), .B(n472), .ZN(n492) );
  NAND2_X1 U584 ( .A1(G214), .A2(n487), .ZN(n637) );
  XOR2_X1 U585 ( .A(G122), .B(G104), .Z(n501) );
  XNOR2_X1 U586 ( .A(n696), .B(n475), .ZN(n486) );
  XOR2_X1 U587 ( .A(KEYINPUT4), .B(KEYINPUT17), .Z(n477) );
  NAND2_X1 U588 ( .A1(G224), .A2(n710), .ZN(n476) );
  XNOR2_X1 U589 ( .A(n477), .B(n476), .ZN(n481) );
  XOR2_X1 U590 ( .A(KEYINPUT72), .B(KEYINPUT85), .Z(n479) );
  XNOR2_X1 U591 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U592 ( .A(n481), .B(n480), .Z(n484) );
  NAND2_X1 U593 ( .A1(n682), .A2(n600), .ZN(n489) );
  AND2_X1 U594 ( .A1(G210), .A2(n487), .ZN(n488) );
  NAND2_X1 U595 ( .A1(n567), .A2(n494), .ZN(n615) );
  NAND2_X1 U596 ( .A1(n651), .A2(n650), .ZN(n525) );
  OR2_X1 U597 ( .A1(n384), .A2(n525), .ZN(n662) );
  XNOR2_X1 U598 ( .A(n495), .B(KEYINPUT31), .ZN(n630) );
  NAND2_X1 U599 ( .A1(n615), .A2(n630), .ZN(n523) );
  XNOR2_X1 U600 ( .A(n497), .B(n496), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n501), .B(KEYINPUT11), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U603 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n508) );
  XNOR2_X1 U604 ( .A(KEYINPUT101), .B(G478), .ZN(n521) );
  XOR2_X1 U605 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n512) );
  XNOR2_X1 U606 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n514), .B(n513), .ZN(n519) );
  XOR2_X1 U608 ( .A(G122), .B(KEYINPUT100), .Z(n517) );
  NAND2_X1 U609 ( .A1(G217), .A2(n515), .ZN(n516) );
  XNOR2_X1 U610 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n519), .B(n518), .ZN(n689) );
  NOR2_X1 U612 ( .A1(G902), .A2(n689), .ZN(n520) );
  XOR2_X1 U613 ( .A(n521), .B(n520), .Z(n524) );
  NOR2_X1 U614 ( .A1(n528), .A2(n524), .ZN(n619) );
  INV_X1 U615 ( .A(n619), .ZN(n631) );
  XNOR2_X2 U616 ( .A(n522), .B(KEYINPUT102), .ZN(n625) );
  INV_X1 U617 ( .A(n625), .ZN(n627) );
  NAND2_X1 U618 ( .A1(n631), .A2(n627), .ZN(n558) );
  INV_X1 U619 ( .A(n524), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n527), .A2(n528), .ZN(n574) );
  NOR2_X1 U621 ( .A1(n525), .A2(n550), .ZN(n526) );
  XNOR2_X1 U622 ( .A(n526), .B(KEYINPUT33), .ZN(n673) );
  NOR2_X1 U623 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U624 ( .A(n529), .B(KEYINPUT103), .ZN(n641) );
  INV_X1 U625 ( .A(KEYINPUT22), .ZN(n530) );
  INV_X1 U626 ( .A(n533), .ZN(n548) );
  OR2_X1 U627 ( .A1(n651), .A2(n548), .ZN(n531) );
  NOR2_X1 U628 ( .A1(n539), .A2(n531), .ZN(n532) );
  NAND2_X1 U629 ( .A1(n532), .A2(n384), .ZN(n618) );
  XNOR2_X1 U630 ( .A(n533), .B(KEYINPUT104), .ZN(n655) );
  AND2_X1 U631 ( .A1(n651), .A2(n655), .ZN(n534) );
  NAND2_X1 U632 ( .A1(n534), .A2(n550), .ZN(n535) );
  XOR2_X1 U633 ( .A(KEYINPUT73), .B(n535), .Z(n536) );
  XNOR2_X1 U634 ( .A(KEYINPUT32), .B(KEYINPUT64), .ZN(n537) );
  XNOR2_X1 U635 ( .A(KEYINPUT77), .B(KEYINPUT45), .ZN(n541) );
  OR2_X1 U636 ( .A1(n710), .A2(n542), .ZN(n543) );
  XOR2_X1 U637 ( .A(KEYINPUT105), .B(n543), .Z(n544) );
  NOR2_X1 U638 ( .A1(G900), .A2(n544), .ZN(n546) );
  NOR2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U640 ( .A(KEYINPUT74), .B(n547), .Z(n568) );
  NOR2_X1 U641 ( .A1(n654), .A2(n548), .ZN(n549) );
  NAND2_X1 U642 ( .A1(n568), .A2(n549), .ZN(n559) );
  XNOR2_X1 U643 ( .A(n592), .B(KEYINPUT107), .ZN(n553) );
  NAND2_X1 U644 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n556), .A2(n651), .ZN(n557) );
  INV_X1 U646 ( .A(n558), .ZN(n643) );
  INV_X1 U647 ( .A(KEYINPUT75), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n643), .A2(n575), .ZN(n565) );
  XNOR2_X1 U649 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n560) );
  XNOR2_X1 U650 ( .A(n561), .B(n560), .ZN(n563) );
  NAND2_X1 U651 ( .A1(n564), .A2(n585), .ZN(n579) );
  INV_X1 U652 ( .A(n579), .ZN(n624) );
  NAND2_X1 U653 ( .A1(n565), .A2(n624), .ZN(n566) );
  NAND2_X1 U654 ( .A1(n566), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n569), .A2(n637), .ZN(n571) );
  NAND2_X1 U656 ( .A1(n595), .A2(n586), .ZN(n573) );
  NOR2_X1 U657 ( .A1(n574), .A2(n573), .ZN(n623) );
  NOR2_X1 U658 ( .A1(KEYINPUT47), .A2(n575), .ZN(n576) );
  NOR2_X1 U659 ( .A1(n623), .A2(n576), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n583) );
  NOR2_X1 U661 ( .A1(KEYINPUT47), .A2(n579), .ZN(n580) );
  NOR2_X1 U662 ( .A1(KEYINPUT75), .A2(n580), .ZN(n581) );
  NOR2_X1 U663 ( .A1(n643), .A2(n581), .ZN(n582) );
  NOR2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U666 ( .A1(n641), .A2(n642), .ZN(n584) );
  XOR2_X1 U667 ( .A(KEYINPUT79), .B(KEYINPUT39), .Z(n587) );
  NAND2_X1 U668 ( .A1(n637), .A2(n590), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT43), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n635) );
  NAND2_X1 U672 ( .A1(n596), .A2(n619), .ZN(n634) );
  NOR2_X1 U673 ( .A1(KEYINPUT2), .A2(n599), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n636), .A2(KEYINPUT2), .ZN(n602) );
  INV_X1 U675 ( .A(n600), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X2 U677 ( .A1(n604), .A2(n603), .ZN(n687) );
  NAND2_X1 U678 ( .A1(n687), .A2(G469), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT125), .ZN(G54) );
  NAND2_X1 U680 ( .A1(n687), .A2(G472), .ZN(n609) );
  XOR2_X1 U681 ( .A(n610), .B(G101), .Z(G3) );
  NOR2_X1 U682 ( .A1(n627), .A2(n615), .ZN(n612) );
  XNOR2_X1 U683 ( .A(G104), .B(KEYINPUT109), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(G6) );
  XOR2_X1 U685 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n614) );
  XNOR2_X1 U686 ( .A(G107), .B(KEYINPUT110), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n617) );
  NOR2_X1 U688 ( .A1(n631), .A2(n615), .ZN(n616) );
  XOR2_X1 U689 ( .A(n617), .B(n616), .Z(G9) );
  XNOR2_X1 U690 ( .A(G110), .B(n618), .ZN(G12) );
  XOR2_X1 U691 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n621) );
  NAND2_X1 U692 ( .A1(n624), .A2(n619), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n621), .B(n620), .ZN(n622) );
  XOR2_X1 U694 ( .A(G128), .B(n622), .Z(G30) );
  XOR2_X1 U695 ( .A(G143), .B(n623), .Z(G45) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n626), .B(G146), .ZN(G48) );
  NOR2_X1 U698 ( .A1(n627), .A2(n630), .ZN(n628) );
  XOR2_X1 U699 ( .A(G113), .B(n628), .Z(n629) );
  XNOR2_X1 U700 ( .A(KEYINPUT112), .B(n629), .ZN(G15) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U702 ( .A(G116), .B(KEYINPUT113), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(G18) );
  XNOR2_X1 U704 ( .A(G134), .B(n634), .ZN(G36) );
  XOR2_X1 U705 ( .A(G140), .B(n635), .Z(G42) );
  XOR2_X1 U706 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n681) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U708 ( .A(KEYINPUT117), .B(n639), .Z(n640) );
  NOR2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n646) );
  NOR2_X1 U710 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n644), .B(KEYINPUT118), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U713 ( .A(KEYINPUT119), .B(n647), .Z(n648) );
  NOR2_X1 U714 ( .A1(n673), .A2(n648), .ZN(n649) );
  XOR2_X1 U715 ( .A(KEYINPUT120), .B(n649), .Z(n668) );
  NOR2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U717 ( .A(KEYINPUT115), .B(n652), .Z(n653) );
  XNOR2_X1 U718 ( .A(KEYINPUT50), .B(n653), .ZN(n659) );
  NAND2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U720 ( .A(n656), .B(KEYINPUT49), .ZN(n657) );
  XNOR2_X1 U721 ( .A(KEYINPUT114), .B(n657), .ZN(n658) );
  NOR2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U723 ( .A1(n660), .A2(n384), .ZN(n661) );
  XNOR2_X1 U724 ( .A(n661), .B(KEYINPUT116), .ZN(n663) );
  NAND2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U726 ( .A(KEYINPUT51), .B(n664), .Z(n665) );
  NAND2_X1 U727 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U729 ( .A(KEYINPUT52), .B(n669), .Z(n670) );
  NOR2_X1 U730 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U733 ( .A(n676), .B(KEYINPUT121), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U735 ( .A1(n679), .A2(n710), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n681), .B(n680), .ZN(G75) );
  NAND2_X1 U737 ( .A1(n687), .A2(G210), .ZN(n683) );
  NAND2_X1 U738 ( .A1(n687), .A2(G475), .ZN(n686) );
  NAND2_X1 U739 ( .A1(G478), .A2(n691), .ZN(n688) );
  XNOR2_X1 U740 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U741 ( .A1(n695), .A2(n690), .ZN(G63) );
  NAND2_X1 U742 ( .A1(G217), .A2(n691), .ZN(n692) );
  XNOR2_X1 U743 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U744 ( .A1(n695), .A2(n694), .ZN(G66) );
  XOR2_X1 U745 ( .A(n696), .B(G107), .Z(n697) );
  NAND2_X1 U746 ( .A1(n698), .A2(n697), .ZN(n706) );
  NAND2_X1 U747 ( .A1(G953), .A2(G224), .ZN(n699) );
  XNOR2_X1 U748 ( .A(KEYINPUT61), .B(n699), .ZN(n700) );
  NAND2_X1 U749 ( .A1(n700), .A2(G898), .ZN(n701) );
  XOR2_X1 U750 ( .A(KEYINPUT126), .B(n701), .Z(n704) );
  NOR2_X1 U751 ( .A1(G953), .A2(n349), .ZN(n703) );
  NOR2_X1 U752 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U753 ( .A(n706), .B(n705), .ZN(G69) );
  XOR2_X1 U754 ( .A(n708), .B(n707), .Z(n712) );
  XNOR2_X1 U755 ( .A(n709), .B(n712), .ZN(n711) );
  NAND2_X1 U756 ( .A1(n711), .A2(n710), .ZN(n716) );
  XNOR2_X1 U757 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U758 ( .A1(n713), .A2(G900), .ZN(n714) );
  NAND2_X1 U759 ( .A1(n714), .A2(G953), .ZN(n715) );
  NAND2_X1 U760 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U761 ( .A(KEYINPUT127), .B(n717), .Z(G72) );
  XNOR2_X1 U762 ( .A(G122), .B(n718), .ZN(G24) );
  XOR2_X1 U763 ( .A(n719), .B(G119), .Z(G21) );
  XOR2_X1 U764 ( .A(n720), .B(G125), .Z(n721) );
  XNOR2_X1 U765 ( .A(KEYINPUT37), .B(n721), .ZN(G27) );
  XOR2_X1 U766 ( .A(n722), .B(G131), .Z(G33) );
  XOR2_X1 U767 ( .A(G137), .B(n723), .Z(G39) );
endmodule

