//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT76), .B(G148gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n203), .B1(new_n214), .B2(new_n204), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n207), .B(new_n208), .C1(new_n213), .C2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT29), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220));
  INV_X1    g019(.A(G211gat), .ZN(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G211gat), .B(G218gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n219), .A3(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n218), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n207), .B1(new_n213), .B2(new_n215), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT29), .B1(new_n227), .B2(new_n228), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT76), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G148gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(G141gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n204), .A2(new_n214), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n210), .B1(new_n202), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G155gat), .B(G162gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(G141gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n210), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n214), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT29), .B1(new_n248), .B2(new_n208), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n236), .B1(new_n249), .B2(new_n229), .ZN(new_n250));
  INV_X1    g049(.A(G228gat), .ZN(new_n251));
  INV_X1    g050(.A(G233gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n231), .B(new_n234), .C1(new_n236), .C2(new_n253), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n255), .B2(new_n256), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n258), .B(new_n265), .C1(new_n260), .C2(KEYINPUT83), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n260), .A2(KEYINPUT83), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT84), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n260), .A2(KEYINPUT83), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n260), .A2(KEYINPUT83), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n258), .A2(new_n265), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277));
  AND2_X1   g076(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n279));
  OAI21_X1  g078(.A(G120gat), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G113gat), .B2(G120gat), .ZN(new_n282));
  INV_X1    g081(.A(G127gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(G134gat), .ZN(new_n284));
  INV_X1    g083(.A(G134gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(G127gat), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n282), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n283), .B2(G134gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT70), .B1(new_n285), .B2(G127gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n283), .A3(G134gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n289), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n280), .A2(new_n287), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n248), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n298), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n297), .A3(new_n280), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(new_n232), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT5), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT3), .B1(new_n243), .B2(new_n247), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n216), .A3(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n310), .A2(new_n216), .A3(new_n304), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(new_n304), .B2(new_n232), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n248), .A2(new_n299), .A3(KEYINPUT4), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n317), .A2(new_n318), .A3(new_n307), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n309), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n318), .A3(new_n307), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n312), .B2(new_n314), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n315), .A2(new_n319), .A3(new_n322), .A4(new_n325), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n321), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G1gat), .B(G29gat), .Z(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G57gat), .B(G85gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n319), .A3(new_n325), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT79), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n327), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n309), .B2(new_n320), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT6), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n334), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n324), .B2(new_n308), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n337), .B2(new_n327), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n345), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n277), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT80), .B1(new_n345), .B2(KEYINPUT6), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n340), .A2(new_n341), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT81), .A4(new_n335), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n329), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(G226gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n252), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT26), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n362), .A2(KEYINPUT26), .ZN(new_n366));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI221_X1 g167(.A(new_n363), .B1(new_n364), .B2(new_n365), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT27), .B(G183gat), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(KEYINPUT67), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT67), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n370), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n376), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n369), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT24), .B1(new_n364), .B2(new_n365), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(G183gat), .A3(G190gat), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n385), .A2(new_n387), .B1(new_n364), .B2(new_n365), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G169gat), .ZN(new_n390));
  INV_X1    g189(.A(G176gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT23), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT65), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n362), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n395));
  INV_X1    g194(.A(new_n362), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n393), .A2(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n389), .B1(new_n398), .B2(KEYINPUT66), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n397), .ZN(new_n400));
  AND4_X1   g199(.A1(new_n394), .A2(new_n390), .A3(new_n391), .A4(KEYINPUT23), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n362), .B2(KEYINPUT23), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(KEYINPUT66), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n384), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(KEYINPUT25), .A3(new_n392), .ZN(new_n406));
  INV_X1    g205(.A(new_n375), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n364), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n385), .A2(new_n387), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n382), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n361), .B1(new_n412), .B2(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n379), .A2(new_n381), .ZN(new_n414));
  INV_X1    g213(.A(new_n369), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n388), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n383), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n416), .B1(new_n420), .B2(new_n410), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n360), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n413), .A2(new_n229), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n360), .B1(new_n421), .B2(new_n217), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT74), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n412), .B2(new_n361), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n360), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n358), .B(new_n423), .C1(new_n428), .C2(new_n229), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n355), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n358), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n427), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n229), .B1(new_n435), .B2(new_n413), .ZN(new_n436));
  INV_X1    g235(.A(new_n423), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n355), .B1(new_n438), .B2(new_n429), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n276), .B1(new_n352), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT73), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n421), .A2(new_n299), .ZN(new_n443));
  INV_X1    g242(.A(G227gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n252), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n416), .B(new_n304), .C1(new_n420), .C2(new_n410), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G15gat), .B(G43gat), .Z(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT72), .ZN(new_n451));
  XOR2_X1   g250(.A(G71gat), .B(G99gat), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n443), .A2(new_n446), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT34), .B1(new_n456), .B2(new_n445), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n445), .B1(new_n443), .B2(new_n446), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n447), .A2(KEYINPUT32), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n453), .B1(new_n447), .B2(new_n448), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n458), .A2(new_n459), .ZN(new_n464));
  AOI211_X1 g263(.A(KEYINPUT34), .B(new_n445), .C1(new_n443), .C2(new_n446), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n461), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n461), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n442), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n442), .B(KEYINPUT36), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n441), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n317), .A2(new_n318), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n307), .B1(new_n315), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n306), .A2(new_n307), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT39), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n334), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n479), .A2(KEYINPUT40), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n343), .B1(new_n338), .B2(new_n321), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT40), .B1(new_n479), .B2(new_n481), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n433), .B2(new_n439), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n485), .B(KEYINPUT85), .C1(new_n433), .C2(new_n439), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n329), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n340), .B2(new_n335), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n423), .C1(new_n428), .C2(new_n229), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n413), .A2(new_n230), .A3(new_n422), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT37), .B(new_n495), .C1(new_n428), .C2(new_n230), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n358), .A2(KEYINPUT38), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n498), .A4(new_n429), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n423), .B1(new_n428), .B2(new_n229), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n358), .B1(new_n500), .B2(KEYINPUT37), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n494), .B1(new_n501), .B2(KEYINPUT87), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n503));
  AOI211_X1 g302(.A(new_n503), .B(new_n358), .C1(new_n500), .C2(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT38), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506));
  INV_X1    g305(.A(new_n340), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n351), .B(new_n429), .C1(new_n507), .C2(new_n483), .ZN(new_n508));
  INV_X1    g307(.A(new_n498), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n511), .A3(new_n276), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n474), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n275), .A2(new_n467), .A3(new_n468), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n352), .A2(new_n515), .A3(new_n440), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n438), .A2(new_n429), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n432), .B1(new_n518), .B2(new_n355), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n519), .B2(new_n492), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n351), .B1(new_n507), .B2(new_n483), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n440), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n520), .A2(new_n521), .A3(new_n524), .A4(new_n515), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n513), .A2(new_n514), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n514), .B1(new_n513), .B2(new_n526), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(G1gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT16), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G1gat), .B2(new_n530), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(G8gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(G8gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(KEYINPUT92), .Z(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n541));
  NOR2_X1   g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT14), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OR4_X1    g345(.A1(new_n540), .A2(new_n541), .A3(new_n543), .A4(new_n546), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n543), .A2(KEYINPUT91), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n540), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT17), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n538), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n537), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT94), .Z(new_n556));
  AND2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n558), .A4(new_n559), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n556), .B1(new_n551), .B2(new_n537), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n558), .B(KEYINPUT13), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT12), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT95), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G99gat), .B(G106gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n552), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n551), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  OAI22_X1  g391(.A1(new_n590), .A2(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT96), .ZN(new_n595));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n591), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n589), .B1(new_n588), .B2(new_n593), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G57gat), .B(G64gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G71gat), .B(G78gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n283), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n537), .B1(KEYINPUT21), .B2(new_n610), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  INV_X1    g418(.A(G155gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n587), .B(new_n610), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n587), .A2(new_n630), .A3(new_n611), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G230gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n252), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n629), .B2(new_n636), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n529), .A2(KEYINPUT97), .A3(new_n577), .A4(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n490), .A2(new_n511), .A3(new_n276), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n348), .A2(new_n349), .A3(new_n335), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n491), .B1(new_n650), .B2(new_n277), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n519), .B1(new_n651), .B2(new_n350), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n471), .B(new_n472), .C1(new_n652), .C2(new_n276), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n526), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT89), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n513), .A2(new_n514), .A3(new_n526), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n577), .A4(new_n647), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n352), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  AND4_X1   g463(.A1(KEYINPUT42), .A2(new_n660), .A3(new_n519), .A4(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT98), .B1(new_n660), .B2(new_n519), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n667));
  AOI211_X1 g466(.A(new_n667), .B(new_n440), .C1(new_n648), .C2(new_n659), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n665), .B1(new_n669), .B2(G8gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n664), .B1(new_n666), .B2(new_n668), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n671), .A2(KEYINPUT99), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT99), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(G1325gat));
  INV_X1    g474(.A(new_n660), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n473), .B(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n467), .A2(new_n468), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n660), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n660), .A2(new_n275), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n689), .B(new_n691), .ZN(G1327gat));
  OR2_X1    g491(.A1(new_n678), .A2(new_n441), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n526), .B1(new_n693), .B2(new_n649), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n604), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n529), .A2(KEYINPUT44), .A3(new_n604), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n627), .ZN(new_n700));
  INV_X1    g499(.A(new_n646), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n577), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n352), .ZN(new_n705));
  INV_X1    g504(.A(new_n577), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n527), .A2(new_n528), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n605), .A2(new_n627), .A3(new_n646), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n544), .A3(new_n661), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n712), .ZN(G1328gat));
  OAI21_X1  g512(.A(G36gat), .B1(new_n704), .B2(new_n440), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n519), .A2(new_n545), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n709), .A2(KEYINPUT104), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT104), .B1(new_n709), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n718), .B2(KEYINPUT46), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721));
  AOI211_X1 g520(.A(KEYINPUT105), .B(new_n721), .C1(new_n716), .C2(new_n717), .ZN(new_n722));
  OAI221_X1 g521(.A(new_n714), .B1(KEYINPUT46), .B2(new_n718), .C1(new_n720), .C2(new_n722), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n678), .A3(new_n698), .A4(new_n703), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT47), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n728), .A3(new_n682), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n727), .B(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n709), .B2(new_n276), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n275), .A2(G50gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n704), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT48), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n733), .B(new_n737), .C1(new_n704), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n628), .A2(new_n577), .A3(new_n701), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n694), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n661), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n440), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n741), .B2(new_n679), .ZN(new_n750));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n682), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n741), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g553(.A1(new_n742), .A2(new_n275), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g555(.A1(new_n706), .A2(KEYINPUT107), .A3(new_n700), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n577), .B2(new_n627), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n694), .A2(new_n604), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT51), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n694), .A2(new_n763), .A3(new_n604), .A4(new_n760), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n579), .A3(new_n661), .A4(new_n646), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n646), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT108), .Z(new_n768));
  NAND3_X1  g567(.A1(new_n699), .A2(new_n661), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G85gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n766), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  NOR3_X1   g573(.A1(new_n701), .A2(G92gat), .A3(new_n440), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n762), .A2(new_n764), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n768), .A2(new_n697), .A3(new_n519), .A4(new_n698), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(KEYINPUT111), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n763), .A2(KEYINPUT110), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n761), .B(new_n783), .Z(new_n784));
  AOI22_X1  g583(.A1(new_n784), .A2(new_n775), .B1(G92gat), .B2(new_n779), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n781), .A2(new_n782), .B1(new_n777), .B2(new_n785), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n699), .A2(new_n678), .A3(new_n768), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G99gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n701), .A2(G99gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n682), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1338gat));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n699), .A2(new_n275), .A3(new_n768), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT112), .B(G106gat), .Z(new_n794));
  NOR3_X1   g593(.A1(new_n701), .A2(G106gat), .A3(new_n276), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n793), .A2(new_n794), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n765), .A2(new_n795), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n792), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n792), .A2(new_n796), .B1(new_n797), .B2(new_n799), .ZN(G1339gat));
  NAND2_X1  g599(.A1(new_n647), .A2(new_n706), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n633), .A2(new_n636), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n635), .B1(new_n631), .B2(new_n632), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n642), .B1(new_n637), .B2(KEYINPUT54), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT113), .B(new_n642), .C1(new_n637), .C2(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n643), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n810), .ZN(new_n814));
  INV_X1    g613(.A(new_n806), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n564), .A2(new_n565), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT115), .Z(new_n824));
  AOI21_X1  g623(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n572), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n576), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n605), .B1(new_n827), .B2(KEYINPUT116), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n822), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n827), .A2(new_n701), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n822), .B2(new_n577), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(new_n604), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n802), .B1(new_n833), .B2(new_n700), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n275), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n352), .A2(new_n519), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n682), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n706), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n834), .A2(new_n352), .ZN(new_n840));
  INV_X1    g639(.A(new_n515), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n519), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n706), .A2(new_n279), .A3(new_n278), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  NOR3_X1   g644(.A1(new_n838), .A2(new_n296), .A3(new_n701), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n646), .A3(new_n842), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n296), .B2(new_n847), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n838), .B2(new_n700), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n627), .A2(new_n283), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n849), .B(KEYINPUT117), .C1(new_n843), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1342gat));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n605), .A2(G134gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n856), .A3(new_n842), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT118), .Z(new_n859));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n842), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n838), .B2(new_n605), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n679), .A2(new_n836), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n834), .B2(new_n276), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n818), .A2(new_n812), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n818), .A2(new_n812), .A3(KEYINPUT119), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n577), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n831), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n604), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n822), .A2(new_n828), .A3(new_n829), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n700), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n801), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n276), .A2(new_n865), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n864), .B1(new_n866), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n209), .B1(new_n879), .B2(new_n577), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n679), .A2(new_n275), .A3(new_n440), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n834), .A2(new_n352), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n209), .A3(new_n577), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT58), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n864), .ZN(new_n886));
  INV_X1    g685(.A(new_n821), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n820), .B1(new_n816), .B2(new_n817), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n577), .B(new_n812), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n604), .B1(new_n889), .B2(new_n872), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n700), .B1(new_n874), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n801), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n275), .ZN(new_n893));
  INV_X1    g692(.A(new_n877), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n875), .B2(new_n801), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n886), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n706), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n883), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n885), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n834), .A2(new_n352), .A3(new_n701), .A4(new_n881), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n212), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n701), .A2(KEYINPUT59), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n886), .B(new_n905), .C1(new_n893), .C2(new_n895), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n903), .A2(new_n237), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n801), .B(KEYINPUT120), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n276), .B1(new_n875), .B2(new_n910), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n911), .A2(KEYINPUT57), .B1(new_n834), .B2(new_n894), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n864), .A2(new_n701), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n901), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n908), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n917), .A2(KEYINPUT121), .A3(new_n904), .A4(new_n906), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(G1345gat));
  OAI21_X1  g718(.A(G155gat), .B1(new_n896), .B2(new_n700), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n882), .A2(new_n620), .A3(new_n627), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  NAND2_X1  g721(.A1(new_n882), .A2(new_n604), .ZN(new_n923));
  INV_X1    g722(.A(G162gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n605), .A2(new_n924), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n896), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n925), .B(new_n930), .C1(new_n896), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n834), .A2(new_n661), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n841), .A2(new_n440), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n577), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n352), .A2(new_n519), .A3(new_n682), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n835), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n390), .A3(new_n706), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n936), .A2(new_n939), .ZN(G1348gat));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n391), .A3(new_n646), .ZN(new_n941));
  OAI21_X1  g740(.A(G176gat), .B1(new_n938), .B2(new_n701), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n627), .A2(new_n371), .A3(new_n378), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n933), .A2(new_n944), .A3(new_n934), .A4(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n892), .A2(new_n276), .A3(new_n627), .A4(new_n937), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G183gat), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n892), .A2(new_n352), .A3(new_n934), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n953), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(G1350gat));
  NAND3_X1  g756(.A1(new_n935), .A2(new_n407), .A3(new_n604), .ZN(new_n958));
  OAI21_X1  g757(.A(G190gat), .B1(new_n938), .B2(new_n605), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n679), .A2(new_n275), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n440), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n933), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g764(.A(KEYINPUT125), .B(G197gat), .Z(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n577), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n678), .A2(new_n661), .A3(new_n440), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n912), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n969), .A2(new_n706), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(new_n966), .ZN(G1352gat));
  OAI21_X1  g770(.A(KEYINPUT127), .B1(new_n969), .B2(new_n701), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n912), .A2(new_n973), .A3(new_n646), .A4(new_n968), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n972), .A2(G204gat), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n701), .A2(G204gat), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n933), .A2(new_n976), .A3(new_n964), .A4(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n892), .A2(new_n352), .A3(new_n964), .A4(new_n977), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT62), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT62), .B1(new_n978), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n975), .A2(new_n983), .ZN(G1353gat));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n221), .A3(new_n627), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n912), .A2(new_n627), .A3(new_n968), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n969), .B2(new_n605), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n965), .A2(new_n222), .A3(new_n604), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


