//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT65), .A2(G134), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n195), .A4(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT0), .B(G128), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(KEYINPUT64), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(G137), .B1(new_n190), .B2(new_n193), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n191), .A2(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n202), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(G131), .C1(new_n217), .C2(new_n218), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n209), .A2(KEYINPUT1), .A3(G146), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n211), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n208), .A3(new_n210), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT69), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n231), .A3(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT30), .B(new_n216), .C1(new_n223), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT2), .A2(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT2), .A3(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(KEYINPUT2), .A2(G113), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n240), .B2(new_n241), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(new_n242), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n209), .A2(KEYINPUT1), .A3(G146), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n204), .B2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n228), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n220), .B2(new_n222), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n206), .A2(new_n214), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n202), .B2(new_n199), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n252), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n234), .A2(new_n251), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n245), .A2(new_n250), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n216), .C1(new_n223), .C2(new_n233), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n261), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n261), .A2(KEYINPUT31), .A3(new_n266), .A4(new_n268), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n251), .B1(new_n259), .B2(new_n257), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n266), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n271), .A2(new_n272), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n271), .A2(new_n272), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n289));
  INV_X1    g103(.A(G472), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n261), .A2(new_n268), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n281), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n281), .B1(new_n268), .B2(new_n278), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n277), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n295), .B(new_n281), .C1(new_n268), .C2(new_n278), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT69), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n231), .B1(new_n226), .B2(new_n228), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n220), .A2(new_n222), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n302), .A2(new_n267), .A3(new_n216), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n267), .B1(new_n302), .B2(new_n216), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT71), .B(new_n290), .C1(new_n296), .C2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n279), .A2(new_n266), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n275), .B1(new_n268), .B2(new_n273), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n295), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n266), .B1(new_n261), .B2(new_n268), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n313), .B2(G472), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n285), .B(new_n289), .C1(new_n307), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G221), .A3(G234), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT73), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G137), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G128), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n322), .A2(G128), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(KEYINPUT23), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT24), .B(G110), .Z(new_n327));
  XNOR2_X1  g141(.A(G119), .B(G128), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT16), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n332), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G146), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(G146), .B1(new_n334), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT72), .B(G110), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n326), .A2(new_n340), .B1(new_n327), .B2(new_n328), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n207), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n336), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n321), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n320), .A2(new_n339), .A3(new_n344), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n348), .B2(KEYINPUT74), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n346), .A2(new_n353), .A3(new_n347), .A4(new_n349), .ZN(new_n354));
  INV_X1    g168(.A(G217), .ZN(new_n355));
  INV_X1    g169(.A(G902), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(G234), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n346), .A2(new_n347), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n357), .A2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n359), .B1(new_n358), .B2(new_n362), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n315), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G214), .B1(G237), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G122), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT82), .Z(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G107), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(G107), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  INV_X1    g193(.A(G101), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n380), .A4(new_n372), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n322), .A3(G116), .ZN(new_n385));
  OAI211_X1 g199(.A(G113), .B(new_n385), .C1(new_n247), .C2(new_n384), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n249), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n376), .A2(new_n379), .A3(new_n372), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n380), .B1(new_n388), .B2(KEYINPUT77), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n376), .A2(new_n379), .A3(new_n390), .A4(new_n372), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n389), .A2(new_n391), .B1(KEYINPUT4), .B2(new_n381), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n250), .B(new_n245), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n393), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT81), .B1(new_n399), .B2(new_n251), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n370), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n251), .A3(KEYINPUT81), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n395), .ZN(new_n403));
  INV_X1    g217(.A(new_n370), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(new_n387), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n370), .C1(new_n396), .C2(new_n400), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n215), .A2(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n229), .A2(new_n332), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(G224), .A3(new_n316), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n316), .A2(G224), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n412), .A2(new_n416), .A3(new_n414), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n406), .A2(new_n408), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n370), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n386), .A2(new_n249), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n382), .A2(KEYINPUT85), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n413), .A2(KEYINPUT7), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(KEYINPUT86), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n411), .B1(KEYINPUT86), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(KEYINPUT86), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n409), .B2(new_n410), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n428), .B(new_n430), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n405), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n421), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n421), .A2(new_n436), .A3(new_n438), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n368), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NOR2_X1   g257(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n256), .A2(new_n382), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n255), .B1(new_n254), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT78), .B(new_n253), .C1(new_n204), .C2(G128), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n382), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n203), .B(new_n445), .C1(new_n447), .C2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n199), .A2(new_n202), .ZN(new_n453));
  AOI21_X1  g267(.A(G128), .B1(new_n208), .B2(new_n210), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n448), .B1(new_n454), .B2(new_n224), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n228), .A3(new_n450), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n383), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(new_n457), .B2(new_n446), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n459));
  OAI21_X1  g273(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n215), .B1(new_n392), .B2(new_n393), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n382), .A2(new_n462), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n230), .A2(new_n464), .A3(new_n232), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n461), .A2(new_n463), .A3(new_n453), .A4(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G140), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n316), .A2(G227), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n467), .B(new_n468), .Z(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n460), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n465), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n258), .B1(new_n397), .B2(new_n398), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n203), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n474), .B2(new_n466), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n443), .B(new_n356), .C1(new_n471), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n458), .A2(new_n459), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n444), .B(new_n453), .C1(new_n457), .C2(new_n446), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n469), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n466), .A2(KEYINPUT80), .A3(new_n470), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT80), .B1(new_n466), .B2(new_n470), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n480), .B(G469), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n443), .A2(new_n356), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT9), .B(G234), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n488), .B2(G902), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT76), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT90), .B1(new_n225), .B2(G143), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n209), .A3(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n209), .A2(G128), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n501), .B2(KEYINPUT91), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(KEYINPUT91), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G134), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n497), .B1(G128), .B2(new_n209), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n190), .A2(new_n193), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(G116), .ZN(new_n510));
  INV_X1    g324(.A(G116), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT89), .A3(G122), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n511), .A2(G122), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n378), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n513), .A2(G107), .A3(new_n515), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n504), .B(new_n507), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n520), .B(new_n516), .C1(new_n513), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n521), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n510), .B2(new_n512), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT92), .B1(new_n524), .B2(new_n515), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n529), .A3(G107), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n505), .A2(new_n506), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n518), .B1(new_n507), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n488), .A2(new_n355), .A3(G953), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n519), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n519), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n356), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G478), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI221_X1 g354(.A(new_n356), .B1(KEYINPUT15), .B2(new_n538), .C1(new_n535), .C2(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(G234), .A2(G237), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(G952), .A3(new_n316), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(G902), .A3(G953), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT21), .B(G898), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G475), .A2(G902), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n337), .A2(new_n338), .ZN(new_n551));
  INV_X1    g365(.A(G237), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n316), .A3(G214), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n209), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT17), .A3(G131), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(G131), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n201), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n551), .B(new_n557), .C1(new_n560), .C2(KEYINPUT17), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g376(.A1(KEYINPUT18), .A2(G131), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n331), .A2(new_n333), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G146), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n343), .ZN(new_n567));
  INV_X1    g381(.A(new_n563), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n556), .A2(KEYINPUT87), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT87), .B1(new_n556), .B2(new_n568), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n564), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(G113), .B(G122), .Z(new_n573));
  XOR2_X1   g387(.A(KEYINPUT88), .B(G104), .Z(new_n574));
  XOR2_X1   g388(.A(new_n573), .B(new_n574), .Z(new_n575));
  AND3_X1   g389(.A1(new_n561), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n342), .A2(KEYINPUT19), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n342), .A2(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n207), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n560), .A2(new_n336), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n550), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT20), .ZN(new_n583));
  INV_X1    g397(.A(new_n575), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n567), .B1(new_n556), .B2(new_n568), .ZN(new_n585));
  INV_X1    g399(.A(new_n571), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n569), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n560), .A2(new_n336), .A3(new_n579), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n561), .A2(new_n572), .A3(new_n575), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT20), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n550), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n575), .B1(new_n561), .B2(new_n572), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n356), .B1(new_n576), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n583), .A2(new_n593), .B1(G475), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n540), .A2(new_n541), .A3(new_n549), .A4(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n442), .A2(new_n493), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n366), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n380), .ZN(G3));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n421), .A2(new_n436), .A3(new_n438), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n438), .B1(new_n421), .B2(new_n436), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n367), .B(new_n549), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n538), .A2(new_n356), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n519), .A2(new_n533), .ZN(new_n607));
  INV_X1    g421(.A(new_n534), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n519), .A2(new_n533), .A3(new_n534), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n606), .B1(new_n611), .B2(new_n538), .ZN(new_n612));
  INV_X1    g426(.A(new_n596), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT33), .B1(new_n535), .B2(new_n536), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n615), .A3(new_n610), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(G478), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n602), .B1(new_n605), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n442), .A2(new_n620), .A3(KEYINPUT94), .A4(new_n549), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n282), .B2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n288), .A2(new_n283), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n487), .A2(new_n365), .A3(new_n491), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT34), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND2_X1  g445(.A1(new_n540), .A2(new_n541), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n592), .B1(new_n591), .B2(new_n550), .ZN(new_n633));
  INV_X1    g447(.A(new_n550), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT20), .B(new_n634), .C1(new_n589), .C2(new_n590), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT95), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n583), .A2(new_n637), .A3(new_n593), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n636), .A2(new_n638), .B1(G475), .B2(new_n595), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n442), .A2(new_n549), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n628), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n625), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n320), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(new_n345), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n361), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n646), .B1(new_n358), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n358), .A2(new_n650), .A3(new_n646), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n597), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n645), .A2(new_n653), .A3(new_n442), .A4(new_n493), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NOR2_X1   g471(.A1(new_n652), .A2(new_n651), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n545), .A2(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n543), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n632), .A2(new_n658), .A3(new_n639), .A4(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n315), .A2(new_n442), .A3(new_n493), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(KEYINPUT99), .B(KEYINPUT39), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n660), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n493), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT100), .Z(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n603), .A2(new_n604), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT38), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n281), .B1(new_n303), .B2(new_n304), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(KEYINPUT98), .B(new_n281), .C1(new_n303), .C2(new_n304), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n674), .A2(new_n269), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n676), .B2(G902), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n289), .A2(new_n285), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n596), .B1(new_n540), .B2(new_n541), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n358), .A2(new_n650), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n367), .A3(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n671), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n668), .A2(new_n669), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  OAI21_X1  g500(.A(new_n367), .B1(new_n603), .B2(new_n604), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n612), .A2(new_n613), .A3(new_n617), .A4(new_n660), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n315), .A3(new_n493), .A4(new_n658), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AOI22_X1  g505(.A1(new_n300), .A2(new_n464), .B1(new_n457), .B2(new_n462), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n453), .B1(new_n692), .B2(new_n461), .ZN(new_n693));
  INV_X1    g507(.A(new_n466), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n469), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n460), .A2(new_n466), .A3(new_n470), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n356), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n489), .A3(new_n476), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n315), .A2(new_n365), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT101), .B1(new_n622), .B2(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n315), .A2(new_n365), .A3(new_n701), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n619), .A4(new_n621), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NOR2_X1   g523(.A1(new_n702), .A2(new_n641), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n511), .ZN(G18));
  NAND4_X1  g525(.A1(new_n315), .A2(new_n442), .A3(new_n653), .A4(new_n701), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  AND2_X1   g527(.A1(new_n271), .A2(new_n272), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n266), .B1(new_n305), .B2(new_n279), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n283), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n623), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n358), .A2(new_n362), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n701), .A3(new_n718), .A4(new_n549), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n680), .B(new_n367), .C1(new_n603), .C2(new_n604), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT102), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n442), .A2(new_n722), .A3(new_n680), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n719), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n509), .ZN(G24));
  AND3_X1   g539(.A1(new_n623), .A2(new_n716), .A3(new_n681), .ZN(new_n726));
  INV_X1    g540(.A(new_n688), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n442), .A3(new_n727), .A4(new_n701), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND2_X1  g543(.A1(new_n487), .A2(new_n489), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n730), .A2(new_n603), .A3(new_n604), .A4(new_n368), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n315), .A3(new_n365), .A4(new_n727), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n732), .A2(KEYINPUT103), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n289), .A2(KEYINPUT104), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n285), .A2(KEYINPUT105), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n288), .A2(new_n741), .A3(KEYINPUT32), .A4(new_n283), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n307), .A2(new_n314), .B1(new_n285), .B2(KEYINPUT105), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n718), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT106), .B(new_n718), .C1(new_n743), .C2(new_n744), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n727), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n738), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NOR3_X1   g568(.A1(new_n603), .A2(new_n604), .A3(new_n368), .ZN(new_n755));
  INV_X1    g569(.A(new_n730), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n315), .A2(new_n365), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n640), .A2(new_n660), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  NAND2_X1  g574(.A1(new_n612), .A2(new_n617), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n596), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT43), .Z(new_n764));
  NOR2_X1   g578(.A1(new_n645), .A2(new_n682), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT108), .Z(new_n767));
  INV_X1    g581(.A(new_n755), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT44), .B1(new_n764), .B2(new_n765), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n489), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n443), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n773), .B2(new_n772), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT107), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(new_n485), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n476), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n771), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n770), .A2(new_n665), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  OR2_X1    g598(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n315), .A2(new_n365), .A3(new_n688), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n755), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  XNOR2_X1  g604(.A(new_n763), .B(KEYINPUT43), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n717), .A2(new_n718), .A3(new_n544), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n671), .A2(new_n368), .A3(new_n701), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT50), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n755), .A2(new_n701), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT115), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n764), .A3(new_n544), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n726), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n801), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n699), .A2(new_n476), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n785), .B(new_n786), .C1(new_n491), .C2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n791), .A2(new_n768), .A3(new_n792), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n804), .A2(new_n365), .A3(new_n544), .A4(new_n679), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n596), .A3(new_n761), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT117), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n809), .A2(new_n810), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n799), .A2(KEYINPUT51), .A3(new_n806), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n805), .A2(new_n749), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT118), .A3(KEYINPUT48), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n316), .A2(G952), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n687), .A2(new_n700), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n793), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n825), .B(new_n828), .C1(new_n824), .C2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n814), .A2(new_n815), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n620), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n819), .A2(new_n820), .A3(new_n823), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n315), .A2(new_n493), .A3(new_n658), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n442), .A2(new_n727), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n662), .B(new_n728), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n681), .B1(new_n543), .B2(new_n659), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n678), .A2(new_n756), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n723), .B2(new_n721), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT52), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n662), .A2(new_n728), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n678), .A2(new_n756), .A3(new_n838), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n722), .B1(new_n442), .B2(new_n680), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n720), .A2(KEYINPUT102), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n842), .A2(new_n843), .A3(new_n690), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n841), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n841), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n605), .A2(KEYINPUT110), .A3(new_n618), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT110), .B1(new_n605), .B2(new_n618), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n853), .A2(new_n627), .A3(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n702), .A2(new_n641), .B1(new_n366), .B2(new_n599), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n540), .A2(new_n541), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n613), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n627), .A2(new_n442), .A3(new_n549), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n712), .A3(new_n654), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n855), .A2(new_n856), .A3(new_n860), .A4(new_n724), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n639), .A3(new_n660), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT111), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n835), .A3(new_n768), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n731), .A2(new_n727), .A3(new_n726), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n757), .B2(new_n758), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n753), .A2(new_n861), .A3(new_n707), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n834), .B1(new_n852), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n732), .A2(KEYINPUT103), .A3(new_n733), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT103), .B1(new_n732), .B2(new_n733), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n867), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n856), .A2(new_n860), .A3(new_n724), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n853), .A2(new_n627), .A3(new_n854), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n707), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n662), .A2(new_n728), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n841), .A2(new_n848), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n878), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n869), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n875), .A2(new_n707), .A3(new_n876), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n862), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n755), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n759), .B(new_n865), .C1(new_n835), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n738), .B2(new_n752), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n886), .A2(new_n891), .A3(new_n881), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT112), .B1(new_n892), .B2(KEYINPUT53), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n878), .A2(new_n881), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n834), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n841), .A2(new_n848), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT113), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n841), .A2(new_n848), .A3(new_n849), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n878), .A2(new_n900), .A3(KEYINPUT53), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n893), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n885), .B1(new_n902), .B2(KEYINPUT54), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n823), .A2(new_n832), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT119), .B1(new_n904), .B2(new_n818), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n833), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(G952), .B2(G953), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n718), .A2(new_n367), .A3(new_n491), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n908), .B(new_n763), .C1(KEYINPUT49), .C2(new_n808), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT109), .Z(new_n911));
  NAND4_X1  g725(.A1(new_n909), .A2(new_n911), .A3(new_n671), .A4(new_n679), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n907), .A2(new_n912), .ZN(G75));
  AOI21_X1  g727(.A(KEYINPUT53), .B1(new_n878), .B2(new_n900), .ZN(new_n914));
  AND4_X1   g728(.A1(KEYINPUT53), .A2(new_n886), .A3(new_n891), .A4(new_n881), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n356), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G210), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n406), .A2(new_n408), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(new_n420), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT56), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n918), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n918), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n316), .A2(G952), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G51));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n914), .B2(new_n915), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n884), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n916), .A2(new_n931), .A3(new_n883), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n485), .B(KEYINPUT57), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n697), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n917), .A2(new_n776), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n927), .B1(new_n935), .B2(new_n936), .ZN(G54));
  NAND2_X1  g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n917), .A2(new_n591), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n591), .B1(new_n917), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n927), .ZN(G60));
  NAND2_X1  g756(.A1(new_n614), .A2(new_n616), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n606), .B(KEYINPUT59), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n930), .A2(new_n932), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n930), .A2(new_n932), .A3(new_n949), .A4(new_n946), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n944), .B1(new_n903), .B2(new_n945), .ZN(new_n952));
  INV_X1    g766(.A(new_n927), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT124), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n948), .A2(new_n950), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n953), .A4(new_n952), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(new_n869), .A2(new_n882), .ZN(new_n960));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT60), .Z(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n953), .B1(new_n963), .B2(new_n360), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n649), .B2(new_n963), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g780(.A1(new_n877), .A2(new_n316), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT125), .Z(new_n968));
  INV_X1    g782(.A(G224), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n547), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n919), .B1(G898), .B2(new_n316), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  AND2_X1   g787(.A1(new_n783), .A2(new_n789), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n723), .A2(new_n721), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n782), .A2(new_n665), .A3(new_n975), .A4(new_n749), .ZN(new_n976));
  INV_X1    g790(.A(new_n837), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n753), .A2(new_n759), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n974), .A2(new_n316), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(G900), .A2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(G227), .A2(G900), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n234), .A2(new_n260), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  NOR2_X1   g798(.A1(new_n577), .A2(new_n578), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AND4_X1   g800(.A1(G953), .A2(new_n981), .A3(new_n982), .A4(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n986), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n979), .B2(new_n980), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n316), .B1(G227), .B2(G900), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n685), .A2(new_n977), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT62), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n755), .B1(new_n858), .B2(new_n620), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n667), .A2(new_n366), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI211_X1 g809(.A(G953), .B(new_n986), .C1(new_n974), .C2(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n989), .A2(new_n990), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n987), .A2(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  NAND3_X1  g814(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n877), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n291), .A2(new_n266), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n927), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n995), .A2(new_n783), .A3(new_n789), .A4(new_n886), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1000), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT127), .B1(new_n1005), .B2(new_n1000), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n266), .B(new_n291), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n292), .A2(new_n269), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n902), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1004), .A2(new_n1008), .A3(new_n1010), .ZN(G57));
endmodule


