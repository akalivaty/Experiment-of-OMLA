//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT2), .B(G113), .Z(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(G116), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT5), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n192), .B2(new_n193), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n191), .A3(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT75), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G104), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n207), .A2(new_n201), .A3(KEYINPUT75), .A4(G104), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n211), .B2(new_n204), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n200), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n202), .A2(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n217));
  AOI211_X1 g031(.A(new_n216), .B(new_n206), .C1(new_n217), .C2(new_n208), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n203), .A2(new_n208), .A3(new_n205), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT76), .B1(new_n219), .B2(G101), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n206), .B1(new_n217), .B2(new_n208), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n189), .A2(new_n194), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(new_n195), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n214), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT80), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT6), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n227), .ZN(new_n230));
  AOI211_X1 g044(.A(new_n230), .B(new_n214), .C1(new_n221), .C2(new_n225), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT81), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n214), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n219), .A2(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n216), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(KEYINPUT76), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n222), .A2(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n224), .A2(new_n195), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n233), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n228), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n233), .B(new_n227), .C1(new_n238), .C2(new_n241), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT6), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G143), .B(G146), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT0), .B(G128), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n261), .A2(new_n249), .A3(new_n251), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n250), .B2(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n249), .A2(KEYINPUT66), .A3(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(G128), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n254), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n259), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G224), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n270), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n242), .A2(new_n275), .A3(new_n243), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n232), .A2(new_n247), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n254), .A2(new_n261), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G125), .ZN(new_n282));
  OAI221_X1 g096(.A(new_n278), .B1(KEYINPUT82), .B2(new_n272), .C1(new_n282), .C2(new_n259), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT7), .B(new_n273), .C1(new_n270), .C2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n227), .B(KEYINPUT8), .Z(new_n287));
  NAND2_X1  g101(.A1(new_n200), .A2(new_n213), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n233), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n231), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n277), .A2(new_n291), .A3(new_n293), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n188), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G475), .A2(G902), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n298), .B(KEYINPUT84), .Z(new_n299));
  INV_X1    g113(.A(KEYINPUT16), .ZN(new_n300));
  INV_X1    g114(.A(G140), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(G125), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n301), .A2(KEYINPUT71), .A3(G125), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(KEYINPUT71), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n304), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n248), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n304), .B(G146), .C1(new_n300), .C2(new_n307), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G214), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n250), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT17), .A3(G131), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(G131), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT17), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n313), .A2(new_n319), .A3(new_n314), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n309), .A2(new_n310), .A3(new_n316), .A4(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G113), .B(G122), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(new_n210), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n307), .A2(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n306), .A2(new_n248), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT18), .A2(G131), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n313), .A2(new_n314), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n315), .A2(KEYINPUT83), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT83), .B1(new_n315), .B2(new_n330), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n327), .B(new_n329), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n322), .A2(new_n324), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT19), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n307), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n306), .A2(KEYINPUT19), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n248), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n317), .A2(new_n320), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n310), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n324), .B1(new_n340), .B2(new_n333), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n299), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n333), .ZN(new_n344));
  INV_X1    g158(.A(new_n324), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n322), .A2(new_n324), .A3(new_n333), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n348), .B2(KEYINPUT20), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT20), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n343), .A3(new_n351), .A4(new_n299), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n324), .B1(new_n322), .B2(new_n333), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n334), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G475), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G952), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(G234), .B2(G237), .ZN(new_n361));
  INV_X1    g175(.A(G234), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  OAI211_X1 g177(.A(G902), .B(G953), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT88), .Z(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT21), .B(G898), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G478), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n369), .A2(KEYINPUT15), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n190), .B2(G122), .ZN(new_n373));
  INV_X1    g187(.A(G122), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT86), .A3(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n190), .A2(G122), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n201), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n201), .B1(new_n376), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n380), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT87), .A3(new_n378), .ZN(new_n383));
  XNOR2_X1  g197(.A(G128), .B(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT13), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n260), .A2(KEYINPUT13), .A3(G143), .ZN(new_n386));
  INV_X1    g200(.A(G134), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n385), .A2(new_n388), .B1(new_n387), .B2(new_n384), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n377), .B(KEYINPUT14), .ZN(new_n391));
  INV_X1    g205(.A(new_n376), .ZN(new_n392));
  OAI21_X1  g206(.A(G107), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n384), .B(new_n387), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n378), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT9), .B(G234), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n397), .A2(new_n398), .A3(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n395), .A3(new_n399), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n370), .B1(new_n403), .B2(new_n354), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n390), .A2(new_n395), .A3(new_n399), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n399), .B1(new_n390), .B2(new_n395), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n354), .B(new_n370), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n358), .A2(new_n368), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G221), .B1(new_n397), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n359), .A2(G227), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT74), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n263), .A2(G128), .B1(new_n249), .B2(new_n251), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(new_n262), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n213), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n260), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n280), .B1(new_n422), .B2(new_n254), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(KEYINPUT77), .A3(new_n209), .A4(new_n212), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n269), .A2(new_n213), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n387), .B2(G137), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n387), .A2(G137), .ZN(new_n430));
  INV_X1    g244(.A(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT11), .A3(G134), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n429), .A2(new_n432), .A3(new_n319), .A4(new_n430), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT12), .B1(new_n436), .B2(KEYINPUT78), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n427), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n421), .A2(new_n424), .B1(new_n269), .B2(new_n213), .ZN(new_n440));
  INV_X1    g254(.A(new_n436), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT10), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n425), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n213), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n256), .B1(new_n222), .B2(new_n223), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n221), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n445), .A2(new_n441), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n417), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n448), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n447), .B1(new_n238), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT10), .B1(new_n421), .B2(new_n424), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n436), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n416), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n455), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n354), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G469), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n450), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n416), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n443), .A2(new_n450), .A3(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT79), .B(G469), .Z(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n354), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n413), .B1(new_n459), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n297), .A2(new_n411), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT73), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n436), .A2(new_n257), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n431), .B2(G134), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT64), .B1(new_n387), .B2(G137), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n431), .A3(G134), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n387), .A2(KEYINPUT65), .A3(G137), .ZN(new_n476));
  AND4_X1   g290(.A1(new_n472), .A2(new_n473), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n435), .B1(new_n477), .B2(new_n319), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n269), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n470), .B(KEYINPUT30), .C1(new_n269), .C2(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n240), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n363), .A2(new_n359), .A3(G210), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT27), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT26), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n484), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT26), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n486), .A2(new_n490), .A3(G101), .ZN(new_n491));
  AOI21_X1  g305(.A(G101), .B1(new_n486), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n240), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n470), .C1(new_n269), .C2(new_n478), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n483), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT31), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n483), .A2(new_n493), .A3(new_n498), .A4(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT67), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n491), .B2(new_n492), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n486), .A2(new_n490), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n206), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n486), .A2(new_n490), .A3(G101), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(KEYINPUT67), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n479), .A2(new_n240), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n495), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n497), .A2(new_n499), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G472), .A2(G902), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n497), .A2(new_n512), .A3(KEYINPUT68), .A4(new_n499), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT69), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n515), .A2(new_n521), .A3(new_n516), .A4(new_n517), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n515), .A2(KEYINPUT32), .A3(new_n516), .A4(new_n517), .ZN(new_n524));
  INV_X1    g338(.A(new_n511), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n501), .A2(new_n505), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n508), .A4(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT29), .B1(new_n511), .B2(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n483), .A2(new_n495), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n493), .B1(new_n531), .B2(new_n526), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n354), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n524), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n523), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G217), .B1(new_n362), .B2(G902), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n309), .A2(new_n310), .ZN(new_n538));
  XOR2_X1   g352(.A(G119), .B(G128), .Z(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT24), .B(G110), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n191), .A2(G128), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT70), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT23), .B1(new_n260), .B2(G119), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(KEYINPUT70), .B2(KEYINPUT23), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(new_n547), .B2(G110), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n539), .A2(new_n540), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n547), .B2(G110), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n310), .A3(new_n326), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT22), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(G137), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(new_n552), .A3(new_n556), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n354), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n537), .B1(new_n560), .B2(KEYINPUT25), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(KEYINPUT25), .B2(new_n560), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n558), .A2(new_n559), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n362), .B2(G217), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n469), .B1(new_n536), .B2(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(KEYINPUT73), .B(new_n566), .C1(new_n523), .C2(new_n535), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n468), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT89), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n206), .ZN(G3));
  NAND3_X1  g386(.A1(new_n515), .A2(new_n354), .A3(new_n517), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G472), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n519), .A2(new_n574), .A3(new_n522), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n466), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n577));
  OR3_X1    g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n575), .B2(new_n576), .ZN(new_n579));
  INV_X1    g393(.A(new_n368), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n297), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n403), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT33), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n403), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n369), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n369), .B1(new_n582), .B2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n358), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n578), .A2(new_n579), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT34), .B(G104), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  XNOR2_X1  g408(.A(new_n342), .B(KEYINPUT20), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n410), .A2(new_n595), .A3(new_n357), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n581), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n578), .A2(new_n579), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  OR2_X1    g414(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(KEYINPUT36), .B2(new_n557), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n564), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n562), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n467), .A2(new_n575), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT37), .B(G110), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  XOR2_X1   g426(.A(KEYINPUT92), .B(G900), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n366), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n361), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n596), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n297), .A2(new_n466), .A3(new_n608), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n536), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G128), .ZN(G30));
  AND3_X1   g435(.A1(new_n277), .A2(new_n291), .A3(new_n293), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n293), .B1(new_n277), .B2(new_n291), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT93), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n295), .A2(new_n625), .A3(new_n296), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT38), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n616), .B(KEYINPUT39), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n466), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n353), .A2(new_n357), .ZN(new_n633));
  NOR4_X1   g447(.A1(new_n608), .A2(new_n633), .A3(new_n188), .A4(new_n409), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n628), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n510), .ZN(new_n636));
  INV_X1    g450(.A(new_n495), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n496), .B1(new_n527), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n354), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n524), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n523), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT94), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G143), .ZN(G45));
  AND3_X1   g460(.A1(new_n358), .A2(new_n589), .A3(new_n616), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n536), .A2(new_n619), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G146), .ZN(G48));
  AOI21_X1  g463(.A(new_n566), .B1(new_n523), .B2(new_n535), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n463), .A2(new_n354), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(KEYINPUT95), .A3(G469), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n654));
  INV_X1    g468(.A(G469), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n412), .A4(new_n465), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT95), .B1(new_n651), .B2(G469), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n654), .A2(new_n653), .A3(new_n655), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n412), .B(new_n465), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT96), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n650), .A2(new_n591), .A3(new_n659), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT41), .B(G113), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  NAND4_X1  g480(.A1(new_n650), .A2(new_n597), .A3(new_n659), .A4(new_n663), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G116), .ZN(G18));
  NAND2_X1  g482(.A1(new_n411), .A2(new_n608), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n523), .B2(new_n535), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n297), .A3(new_n659), .A4(new_n663), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G119), .ZN(G21));
  NAND2_X1  g486(.A1(new_n513), .A2(new_n516), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n574), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n566), .A3(new_n368), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n409), .B1(new_n353), .B2(new_n357), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n676), .B(new_n187), .C1(new_n622), .C2(new_n623), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n297), .A2(KEYINPUT97), .A3(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n675), .A2(new_n681), .A3(new_n659), .A4(new_n663), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G122), .ZN(G24));
  AOI22_X1  g497(.A1(new_n573), .A2(G472), .B1(new_n516), .B2(new_n513), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n684), .A2(new_n608), .A3(new_n647), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n663), .A3(new_n297), .A4(new_n659), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G125), .ZN(G27));
  AND2_X1   g501(.A1(new_n518), .A2(new_n520), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n524), .A2(new_n534), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n567), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT98), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n458), .B2(G469), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n451), .A2(new_n457), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n655), .A2(KEYINPUT98), .A3(G902), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n465), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n622), .A2(new_n623), .A3(new_n188), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n647), .A3(new_n697), .A4(new_n412), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n690), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n696), .A2(new_n412), .A3(new_n697), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n650), .A2(new_n647), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n700), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n319), .ZN(G33));
  NAND3_X1  g518(.A1(new_n650), .A2(new_n618), .A3(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G134), .ZN(G36));
  NAND2_X1  g520(.A1(new_n633), .A2(new_n589), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT43), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n712));
  NAND3_X1  g526(.A1(new_n633), .A2(new_n589), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n714), .A2(new_n608), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n710), .A2(new_n713), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT103), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n575), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n697), .B(KEYINPUT104), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n575), .A4(new_n717), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n455), .A2(new_n450), .A3(new_n456), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n453), .A2(new_n454), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n441), .A2(new_n725), .B1(new_n439), .B2(new_n442), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n724), .B1(new_n726), .B2(new_n417), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n655), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n693), .A2(KEYINPUT99), .A3(KEYINPUT45), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(G469), .A2(G902), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT46), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT100), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n734), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n465), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n412), .A3(new_n629), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT101), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(KEYINPUT101), .A3(new_n412), .A4(new_n629), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n723), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT105), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G137), .ZN(G39));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n740), .A2(new_n748), .A3(new_n412), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n748), .B1(new_n740), .B2(new_n412), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n647), .A2(new_n697), .A3(new_n566), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n536), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT106), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n301), .ZN(G42));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n357), .A2(new_n595), .A3(new_n409), .A4(new_n616), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n697), .A2(new_n466), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n536), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n693), .A2(new_n694), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n655), .B1(new_n727), .B2(new_n354), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n691), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n413), .B1(new_n765), .B2(new_n465), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n647), .A3(new_n684), .A4(new_n697), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n609), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n650), .A2(new_n618), .A3(new_n701), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT110), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n698), .A2(new_n674), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n760), .B1(new_n523), .B2(new_n535), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n608), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n705), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n664), .A2(new_n671), .A3(new_n667), .A4(new_n682), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n703), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n633), .A2(new_n410), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n581), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n578), .A2(new_n579), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n610), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n536), .A2(new_n567), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT73), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n650), .A2(new_n469), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n467), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n578), .A2(new_n579), .A3(new_n591), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT109), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n570), .A2(new_n790), .A3(new_n592), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n783), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n686), .A2(new_n620), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n608), .A2(new_n617), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n696), .A3(new_n412), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n766), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n679), .A2(new_n680), .B1(new_n523), .B2(new_n642), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n686), .A2(KEYINPUT111), .A3(new_n620), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n795), .A2(new_n648), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n803), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n686), .A2(new_n620), .A3(new_n648), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n796), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n779), .A2(new_n792), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n807), .A2(new_n620), .A3(new_n648), .A4(new_n686), .ZN(new_n815));
  INV_X1    g629(.A(new_n809), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n796), .B1(new_n816), .B2(new_n804), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n779), .A2(new_n818), .A3(new_n792), .A4(KEYINPUT53), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n758), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n783), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n570), .A2(new_n790), .A3(new_n592), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n790), .B1(new_n570), .B2(new_n592), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n703), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n664), .A2(new_n671), .A3(new_n667), .A4(new_n682), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT110), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n774), .B1(new_n773), .B2(new_n705), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n824), .A2(new_n829), .A3(new_n817), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT113), .B1(new_n830), .B2(KEYINPUT53), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n779), .A2(new_n792), .A3(KEYINPUT53), .A4(new_n811), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n833), .B(new_n834), .C1(new_n830), .C2(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n663), .A2(new_n659), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n697), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n697), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n644), .A2(new_n567), .A3(new_n361), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n358), .A2(new_n589), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n716), .A2(new_n361), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n567), .B(new_n684), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n628), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n188), .A3(new_n837), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT50), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n852), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n855), .ZN(new_n860));
  AND4_X1   g674(.A1(KEYINPUT50), .A2(new_n857), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n847), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n850), .A2(new_n851), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n842), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n842), .B2(new_n866), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n608), .B(new_n684), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n657), .A2(new_n465), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT107), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n412), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n721), .B(new_n859), .C1(new_n752), .C2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n863), .A2(KEYINPUT51), .A3(new_n869), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n874), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n877), .B2(new_n862), .ZN(new_n878));
  INV_X1    g692(.A(new_n690), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n867), .B2(new_n868), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n360), .B(KEYINPUT118), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n837), .A2(new_n297), .ZN(new_n883));
  OAI221_X1 g697(.A(new_n882), .B1(new_n883), .B2(new_n852), .C1(new_n844), .C2(new_n590), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT119), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n875), .A2(new_n878), .A3(new_n881), .A4(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n836), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n872), .A2(KEYINPUT49), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT108), .Z(new_n889));
  OR4_X1    g703(.A1(new_n566), .A2(new_n707), .A3(new_n188), .A4(new_n413), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n628), .B(new_n890), .C1(new_n872), .C2(KEYINPUT49), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n644), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(G75));
  NAND3_X1  g707(.A1(new_n779), .A2(new_n818), .A3(new_n792), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n813), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n354), .B1(new_n895), .B2(new_n834), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G210), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n232), .A2(new_n247), .A3(new_n276), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n274), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n897), .B2(new_n898), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n359), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n835), .A2(KEYINPUT120), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n895), .A2(new_n907), .A3(new_n833), .A4(new_n834), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n824), .A2(new_n829), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT53), .B1(new_n909), .B2(new_n818), .ZN(new_n910));
  INV_X1    g724(.A(new_n834), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT54), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n734), .B(KEYINPUT57), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n463), .ZN(new_n916));
  INV_X1    g730(.A(new_n896), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(new_n733), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n904), .B1(new_n916), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n347), .A3(new_n346), .ZN(new_n921));
  INV_X1    g735(.A(new_n904), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(new_n350), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G60));
  AND2_X1   g738(.A1(new_n583), .A2(new_n585), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n836), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n925), .A2(new_n927), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n922), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n895), .B2(new_n834), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(new_n563), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n604), .A2(new_n606), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n904), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT121), .B1(new_n935), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n936), .B(new_n938), .C1(new_n940), .C2(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  NAND2_X1  g758(.A1(new_n792), .A2(new_n826), .ZN(new_n945));
  NAND2_X1  g759(.A1(G224), .A2(G953), .ZN(new_n946));
  OAI22_X1  g760(.A1(new_n945), .A2(G953), .B1(new_n367), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n899), .B1(G898), .B2(new_n359), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n947), .B(new_n948), .Z(G69));
  AOI21_X1  g763(.A(new_n359), .B1(G227), .B2(G900), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n481), .A2(new_n482), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT122), .Z(new_n952));
  NOR2_X1   g766(.A1(new_n336), .A2(new_n337), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(G900), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n743), .A2(new_n744), .ZN(new_n956));
  INV_X1    g770(.A(new_n723), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n690), .B1(new_n679), .B2(new_n680), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n648), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n793), .B2(new_n794), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(new_n805), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n703), .A2(new_n769), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n959), .A2(new_n755), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n955), .B1(new_n964), .B2(G953), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(KEYINPUT126), .B(new_n955), .C1(new_n964), .C2(G953), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n954), .B(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n785), .A2(new_n786), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n630), .B1(new_n590), .B2(new_n780), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n971), .A2(new_n697), .A3(new_n972), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n745), .A2(KEYINPUT124), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n645), .A2(new_n805), .A3(new_n961), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT124), .B1(new_n745), .B2(new_n973), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n974), .A2(new_n755), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(new_n359), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n950), .B1(new_n969), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n950), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n982), .B(new_n965), .C1(new_n980), .C2(KEYINPUT125), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n979), .B2(new_n945), .ZN(new_n988));
  INV_X1    g802(.A(new_n493), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n531), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n964), .B2(new_n945), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n531), .A2(new_n989), .ZN(new_n995));
  OAI211_X1 g809(.A(KEYINPUT127), .B(new_n987), .C1(new_n964), .C2(new_n945), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n991), .A2(new_n922), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n820), .A2(new_n831), .ZN(new_n999));
  INV_X1    g813(.A(new_n987), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n999), .A2(new_n995), .A3(new_n990), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n998), .A2(new_n1001), .ZN(G57));
endmodule


