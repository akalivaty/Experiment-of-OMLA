//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1316, new_n1317, new_n1318, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n209), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT64), .B(G77), .Z(new_n222));
  AOI21_X1  g0022(.A(new_n221), .B1(G244), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT65), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n226), .B(new_n227), .C1(new_n223), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n214), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n211), .B(new_n217), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n236), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT67), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1698), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(G222), .A2(new_n255), .B1(new_n222), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(new_n254), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT69), .B(G223), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n208), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(new_n264), .B2(new_n208), .ZN(new_n268));
  AND2_X1   g0068(.A1(G1), .A2(G13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n268), .A2(new_n271), .A3(new_n273), .A4(G274), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n268), .A2(new_n271), .A3(G226), .A4(new_n272), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(G190), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(KEYINPUT73), .B(G200), .Z(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n265), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n259), .B2(new_n262), .ZN(new_n282));
  OAI211_X1 g0082(.A(KEYINPUT74), .B(new_n280), .C1(new_n282), .C2(new_n276), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n209), .A3(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n202), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n208), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G1), .B2(new_n209), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n286), .B1(new_n290), .B2(new_n202), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT8), .ZN(new_n294));
  INV_X1    g0094(.A(G58), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(KEYINPUT70), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT8), .A3(G58), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n298), .A3(new_n209), .A4(G33), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n289), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT9), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n288), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n284), .A2(G1), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n288), .B1(new_n212), .B2(G20), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(G50), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n278), .A2(new_n283), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n266), .A2(new_n277), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT74), .B1(new_n313), .B2(new_n280), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT10), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n282), .A2(new_n276), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(G190), .B1(new_n301), .B2(new_n310), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT74), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n316), .B2(new_n279), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n317), .A2(new_n319), .A3(new_n320), .A4(new_n283), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n313), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n303), .A2(new_n308), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  OAI211_X1 g0131(.A(G232), .B(new_n331), .C1(new_n256), .C2(new_n257), .ZN(new_n332));
  OAI211_X1 g0132(.A(G238), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n253), .A2(G107), .A3(new_n254), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(new_n265), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n268), .A2(new_n271), .A3(G244), .A4(new_n272), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n274), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT71), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n274), .A2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n265), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n280), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G77), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n290), .A2(new_n345), .B1(new_n222), .B2(new_n305), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT8), .B(G58), .Z(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n292), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT64), .B(G77), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n209), .A2(G33), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n348), .B1(new_n209), .B2(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n352), .B2(new_n288), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n336), .A2(KEYINPUT71), .A3(new_n338), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n341), .B1(new_n340), .B2(new_n342), .ZN(new_n356));
  OAI21_X1  g0156(.A(G190), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n339), .A2(new_n343), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT72), .A3(G190), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n354), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n326), .ZN(new_n363));
  INV_X1    g0163(.A(new_n353), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n339), .A2(new_n323), .A3(new_n343), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G226), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n331), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n238), .A2(G1698), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n370), .C1(new_n256), .C2(new_n257), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G97), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n265), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n268), .A2(new_n271), .A3(G238), .A4(new_n272), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n274), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n378), .B1(new_n377), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(G169), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n281), .B1(new_n373), .B2(KEYINPUT75), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n380), .B1(new_n390), .B2(new_n376), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(new_n378), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n378), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n388), .A2(new_n392), .A3(G179), .A4(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n385), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n345), .B2(new_n350), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n288), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT77), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n400), .A3(new_n288), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT11), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT11), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n404), .A3(new_n401), .ZN(new_n405));
  OR3_X1    g0205(.A1(new_n305), .A2(KEYINPUT12), .A3(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT12), .B1(new_n305), .B2(G68), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n406), .A2(new_n407), .B1(G68), .B2(new_n307), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G200), .B1(new_n382), .B2(new_n383), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n388), .A2(new_n392), .A3(G190), .A4(new_n393), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n395), .A2(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT78), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n330), .B(new_n367), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n253), .A2(new_n209), .A3(new_n254), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT7), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n254), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(KEYINPUT79), .A3(new_n418), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(G68), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n295), .A2(new_n219), .ZN(new_n425));
  OAI21_X1  g0225(.A(G20), .B1(new_n425), .B2(new_n201), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n292), .A2(G159), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT16), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n289), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n219), .B1(new_n419), .B2(new_n421), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT80), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT80), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n429), .C1(new_n432), .C2(new_n428), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n296), .A2(new_n298), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n305), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n307), .B2(new_n438), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n268), .A2(G274), .A3(new_n271), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n368), .A2(G1698), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G223), .B2(G1698), .ZN(new_n444));
  INV_X1    g0244(.A(G87), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n444), .A2(new_n258), .B1(new_n252), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n442), .A2(new_n273), .B1(new_n446), .B2(new_n265), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n268), .A2(new_n271), .A3(G232), .A4(new_n272), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(G179), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G223), .A2(G1698), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n368), .B2(G1698), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n260), .B1(G33), .B2(G87), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n448), .B(new_n274), .C1(new_n452), .C2(new_n281), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G169), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(KEYINPUT18), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n437), .A2(new_n440), .B1(new_n454), .B2(new_n449), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT18), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n441), .A2(new_n455), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  INV_X1    g0265(.A(G190), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n447), .A2(new_n465), .A3(new_n466), .A4(new_n448), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT82), .B1(new_n453), .B2(G190), .ZN(new_n468));
  INV_X1    g0268(.A(G200), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n437), .A2(new_n471), .A3(new_n440), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT83), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(KEYINPUT17), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n464), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n395), .A2(new_n409), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n413), .A2(new_n411), .A3(new_n410), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n478), .A2(new_n415), .A3(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n416), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n260), .A2(G244), .A3(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  OAI211_X1 g0284(.A(G238), .B(new_n331), .C1(new_n256), .C2(new_n257), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n265), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n264), .A2(new_n267), .A3(new_n208), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT68), .B1(new_n269), .B2(new_n270), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  OR3_X1    g0291(.A1(new_n491), .A2(G1), .A3(G274), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(G1), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n490), .B(new_n492), .C1(G250), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n280), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n260), .A2(new_n209), .A3(G68), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  INV_X1    g0298(.A(G97), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n350), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n445), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT89), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n445), .A2(new_n499), .A3(new_n502), .A4(KEYINPUT89), .ZN(new_n506));
  NAND3_X1  g0306(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n505), .A2(new_n506), .B1(new_n209), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n288), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n351), .A2(new_n285), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n289), .B(new_n305), .C1(G1), .C2(new_n252), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G87), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n487), .A2(new_n494), .A3(G190), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n496), .A2(new_n511), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n351), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n509), .A3(new_n510), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n487), .A2(new_n494), .A3(new_n326), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n487), .A2(new_n494), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(G169), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n285), .A2(KEYINPUT25), .A3(new_n502), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT25), .B1(new_n285), .B2(new_n502), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n512), .A2(new_n502), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n209), .B2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n502), .A2(KEYINPUT23), .A3(G20), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n209), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n260), .A2(new_n536), .A3(new_n209), .A4(G87), .ZN(new_n537));
  AOI211_X1 g0337(.A(KEYINPUT24), .B(new_n533), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n537), .ZN(new_n540));
  INV_X1    g0340(.A(new_n533), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n288), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT94), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT94), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n288), .C1(new_n538), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n527), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G41), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n212), .B(G45), .C1(new_n548), .C2(KEYINPUT5), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT5), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G41), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n493), .A2(KEYINPUT86), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(KEYINPUT87), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT87), .B1(new_n551), .B2(new_n554), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n548), .A2(KEYINPUT5), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n268), .A2(new_n271), .A3(G274), .A4(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(new_n558), .A3(new_n554), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n490), .A3(G264), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n563));
  OAI211_X1 g0363(.A(G250), .B(new_n331), .C1(new_n256), .C2(new_n257), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G294), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n265), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n469), .B1(new_n560), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT95), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT95), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n571), .B(new_n469), .C1(new_n560), .C2(new_n568), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n562), .A2(new_n567), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT87), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n549), .A2(new_n550), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT86), .B1(new_n493), .B2(new_n553), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(new_n442), .A3(new_n558), .A4(new_n555), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n466), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n523), .B1(new_n547), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n499), .A2(new_n502), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G97), .A2(G107), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(KEYINPUT6), .A2(G97), .ZN(new_n586));
  OR3_X1    g0386(.A1(new_n586), .A2(KEYINPUT84), .A3(G107), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT84), .B1(new_n586), .B2(G107), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n419), .A2(new_n421), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(KEYINPUT85), .A3(G107), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n502), .B1(new_n419), .B2(new_n421), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(KEYINPUT85), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n288), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n305), .A2(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n513), .B2(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G244), .B(new_n331), .C1(new_n256), .C2(new_n257), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT4), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n331), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G283), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n265), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n561), .A2(new_n490), .A3(G257), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n578), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n323), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n607), .A2(new_n578), .A3(new_n608), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n326), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n599), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n607), .A2(new_n608), .A3(new_n578), .A4(new_n466), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n611), .B2(G200), .ZN(new_n615));
  INV_X1    g0415(.A(new_n598), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n594), .A2(KEYINPUT85), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n592), .A3(new_n590), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n618), .B2(new_n288), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT88), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n615), .A2(KEYINPUT88), .A3(new_n619), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n581), .B(new_n613), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n527), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n540), .A2(new_n541), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT24), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n540), .A2(new_n539), .A3(new_n541), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n545), .B1(new_n627), .B2(new_n288), .ZN(new_n628));
  INV_X1    g0428(.A(new_n546), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n573), .A2(new_n578), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n323), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n573), .A2(new_n326), .A3(new_n578), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n561), .A2(new_n490), .A3(G270), .ZN(new_n637));
  OAI211_X1 g0437(.A(G264), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n638));
  OAI211_X1 g0438(.A(G257), .B(new_n331), .C1(new_n256), .C2(new_n257), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n253), .A2(G303), .A3(new_n254), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n265), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(G200), .B1(new_n560), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n578), .A2(G190), .A3(new_n637), .A4(new_n642), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G116), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n287), .A2(new_n208), .B1(G20), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(G20), .B1(G33), .B2(G283), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n252), .A2(G97), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  OAI211_X1 g0453(.A(KEYINPUT20), .B(new_n648), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT91), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n649), .A2(new_n650), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT90), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(KEYINPUT91), .A3(KEYINPUT20), .A4(new_n648), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT20), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n656), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n305), .A2(new_n647), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n513), .B2(new_n647), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT93), .B1(new_n646), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n665), .A2(new_n667), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT93), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n645), .A4(new_n644), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT21), .ZN(new_n674));
  OAI21_X1  g0474(.A(G169), .B1(new_n560), .B2(new_n643), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n637), .A2(new_n642), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n323), .B1(new_n677), .B2(new_n578), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT21), .B1(new_n678), .B2(new_n668), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(G179), .A3(new_n578), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT92), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  AND4_X1   g0482(.A1(G179), .A2(new_n578), .A3(new_n637), .A4(new_n642), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n668), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n636), .A2(new_n673), .A3(new_n680), .A4(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n482), .A2(new_n622), .A3(new_n687), .ZN(G372));
  INV_X1    g0488(.A(new_n328), .ZN(new_n689));
  INV_X1    g0489(.A(new_n322), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n463), .A2(new_n456), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n395), .A2(new_n409), .B1(new_n479), .B2(new_n366), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n476), .B1(new_n692), .B2(KEYINPUT96), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n479), .A2(new_n366), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n478), .A2(KEYINPUT96), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n691), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT97), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n690), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(KEYINPUT97), .B(new_n691), .C1(new_n693), .C2(new_n695), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n522), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n599), .A2(new_n610), .A3(new_n612), .ZN(new_n702));
  INV_X1    g0502(.A(new_n523), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(KEYINPUT26), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT26), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n613), .B2(new_n523), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n674), .B1(new_n670), .B2(new_n675), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n678), .A2(KEYINPUT21), .A3(new_n668), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n683), .A2(new_n668), .A3(new_n684), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n684), .B1(new_n683), .B2(new_n668), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n708), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n544), .A2(new_n546), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n634), .B1(new_n713), .B2(new_n623), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n707), .B1(new_n622), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n481), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n700), .A2(new_n717), .ZN(G369));
  INV_X1    g0518(.A(KEYINPUT98), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n304), .A2(new_n209), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(G213), .ZN(new_n723));
  INV_X1    g0523(.A(G343), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n668), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n673), .A2(new_n680), .A3(new_n686), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n712), .A2(new_n668), .A3(new_n725), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n719), .B1(new_n729), .B2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  AOI211_X1 g0531(.A(KEYINPUT98), .B(new_n731), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n630), .A2(new_n725), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n547), .A2(new_n580), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n636), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n714), .A2(new_n725), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n725), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n714), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n712), .A2(new_n741), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n740), .A2(new_n745), .ZN(G399));
  INV_X1    g0546(.A(new_n215), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G41), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n505), .A2(new_n647), .A3(new_n506), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n749), .A2(G1), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n206), .B2(new_n749), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n677), .A2(new_n578), .ZN(new_n755));
  AOI21_X1  g0555(.A(G179), .B1(new_n487), .B2(new_n494), .ZN(new_n756));
  AND4_X1   g0556(.A1(new_n609), .A2(new_n631), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n609), .A2(new_n568), .A3(new_n495), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT99), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n683), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n681), .A2(KEYINPUT99), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT30), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n758), .A2(new_n760), .A3(new_n761), .A4(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n741), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n669), .A2(new_n672), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n767), .A2(new_n712), .A3(new_n714), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n615), .A2(new_n619), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT88), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n615), .A2(KEYINPUT88), .A3(new_n619), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n702), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n768), .A2(new_n773), .A3(new_n581), .A4(new_n741), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n766), .B1(new_n774), .B2(KEYINPUT31), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(KEYINPUT31), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(G330), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n636), .A2(new_n686), .A3(new_n680), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n773), .A2(new_n780), .A3(new_n581), .ZN(new_n781));
  AOI211_X1 g0581(.A(KEYINPUT29), .B(new_n725), .C1(new_n781), .C2(new_n707), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT29), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n716), .B2(new_n741), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n754), .B1(new_n787), .B2(G1), .ZN(G364));
  NOR2_X1   g0588(.A1(new_n284), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n212), .B1(new_n789), .B2(G45), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n748), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n733), .B(new_n793), .C1(G330), .C2(new_n729), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n215), .A2(new_n260), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n795), .A2(new_n796), .B1(G116), .B2(new_n215), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n249), .A2(G45), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n747), .A2(new_n260), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n491), .B2(new_n207), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n208), .B1(G20), .B2(new_n323), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n792), .B1(new_n803), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(G20), .A2(G179), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT102), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G190), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G200), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n466), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n469), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G58), .A2(new_n818), .B1(new_n820), .B2(G68), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n817), .A2(new_n469), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n819), .A2(G200), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G50), .A2(new_n822), .B1(new_n823), .B2(new_n222), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n466), .A2(G179), .A3(G200), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n209), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n260), .B1(new_n826), .B2(new_n499), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n209), .A2(G179), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n280), .A2(G190), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n827), .B1(new_n830), .B2(G87), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n280), .A2(new_n466), .A3(new_n828), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR4_X1   g0633(.A1(new_n209), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n834), .A2(KEYINPUT32), .A3(G159), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT32), .ZN(new_n836));
  INV_X1    g0636(.A(new_n834), .ZN(new_n837));
  INV_X1    g0637(.A(G159), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n833), .A2(G107), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n821), .A2(new_n824), .A3(new_n831), .A4(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n826), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(G294), .B1(G329), .B2(new_n834), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  INV_X1    g0644(.A(new_n823), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n843), .B1(new_n844), .B2(new_n832), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G326), .B2(new_n822), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n260), .B1(new_n830), .B2(G303), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT103), .Z(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(KEYINPUT33), .B(G317), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G322), .A2(new_n818), .B1(new_n820), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT104), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n814), .B1(new_n855), .B2(new_n808), .ZN(new_n856));
  INV_X1    g0656(.A(new_n811), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n729), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n794), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G396));
  NAND2_X1  g0660(.A1(new_n716), .A2(new_n741), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n353), .A2(new_n741), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n362), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n725), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n725), .B(new_n868), .C1(new_n781), .C2(new_n707), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n779), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT105), .Z(new_n874));
  OAI211_X1 g0674(.A(new_n874), .B(new_n793), .C1(new_n779), .C2(new_n872), .ZN(new_n875));
  INV_X1    g0675(.A(new_n808), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n810), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n792), .B1(new_n877), .B2(G77), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n818), .B1(new_n823), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(new_n822), .ZN(new_n881));
  INV_X1    g0681(.A(G150), .ZN(new_n882));
  INV_X1    g0682(.A(new_n820), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n879), .B1(new_n880), .B2(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT34), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n830), .A2(G50), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n833), .A2(G68), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n842), .A2(G58), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n258), .B1(new_n834), .B2(G132), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n258), .B1(new_n837), .B2(new_n846), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(G97), .B2(new_n842), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n833), .A2(G87), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n892), .B(new_n893), .C1(new_n502), .C2(new_n829), .ZN(new_n894));
  AOI22_X1  g0694(.A1(G294), .A2(new_n818), .B1(new_n822), .B2(G303), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n895), .B1(new_n647), .B2(new_n845), .C1(new_n844), .C2(new_n883), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n885), .A2(new_n890), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n878), .B1(new_n897), .B2(new_n808), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n810), .B2(new_n869), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n875), .A2(new_n899), .ZN(G384));
  OR2_X1    g0700(.A1(new_n589), .A2(KEYINPUT35), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n589), .A2(KEYINPUT35), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n901), .A2(G116), .A3(new_n210), .A4(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT36), .Z(new_n904));
  OAI211_X1 g0704(.A(new_n222), .B(new_n207), .C1(new_n295), .C2(new_n219), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n202), .A2(G68), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n212), .B(G13), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n476), .A2(new_n691), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n723), .B1(new_n437), .B2(new_n440), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n461), .A2(new_n472), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT106), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n461), .A2(KEYINPUT106), .A3(new_n472), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n723), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n441), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n461), .A2(new_n919), .A3(new_n912), .A4(new_n472), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT107), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n472), .A4(new_n461), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n911), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n424), .A2(new_n430), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n288), .ZN(new_n930));
  INV_X1    g0730(.A(new_n428), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT16), .B1(new_n424), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n440), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n918), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n455), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n472), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT37), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n920), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n464), .A2(new_n476), .ZN(new_n940));
  OAI211_X1 g0740(.A(KEYINPUT38), .B(new_n939), .C1(new_n940), .C2(new_n935), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT39), .B1(new_n928), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n935), .B1(new_n464), .B2(new_n476), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n938), .A2(new_n920), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n927), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n478), .A2(new_n725), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n942), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n409), .A2(new_n725), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n414), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n414), .A2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n871), .B2(new_n866), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n941), .A2(new_n945), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n955), .A2(new_n956), .B1(new_n691), .B2(new_n918), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n481), .B1(new_n782), .B2(new_n784), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n700), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n958), .B(new_n960), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n869), .B1(new_n951), .B2(new_n952), .ZN(new_n962));
  INV_X1    g0762(.A(new_n766), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n622), .A2(new_n687), .A3(new_n725), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT31), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT108), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n766), .A2(new_n967), .A3(KEYINPUT31), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n766), .B2(KEYINPUT31), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n962), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n922), .A2(new_n924), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n437), .A2(new_n471), .A3(new_n440), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n914), .B1(new_n973), .B2(new_n458), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(new_n916), .A3(new_n919), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT37), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n972), .A2(new_n976), .B1(new_n910), .B2(new_n909), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n941), .B1(new_n977), .B2(KEYINPUT38), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT40), .B1(new_n941), .B2(new_n945), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n979), .A2(KEYINPUT40), .B1(new_n971), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n966), .A2(new_n970), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(new_n481), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n731), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n984), .B2(new_n982), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n961), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n212), .B2(new_n789), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n961), .A2(new_n986), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n908), .B1(new_n988), .B2(new_n989), .ZN(G367));
  NOR2_X1   g0790(.A1(new_n737), .A2(new_n743), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n599), .A2(new_n725), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n613), .B(new_n992), .C1(new_n621), .C2(new_n620), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n613), .A2(new_n741), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n613), .B1(new_n993), .B2(new_n636), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n997), .A2(KEYINPUT42), .B1(new_n741), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n511), .A2(new_n514), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n725), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n703), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n522), .B2(new_n1002), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n998), .A2(new_n1000), .B1(KEYINPUT43), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n733), .B1(new_n738), .B2(new_n737), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n996), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1007), .B(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n748), .B(KEYINPUT41), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n729), .A2(G330), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT98), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n725), .B1(new_n680), .B2(new_n686), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1015), .A2(new_n736), .A3(new_n636), .A4(new_n735), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n729), .A2(new_n719), .A3(G330), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1014), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n730), .B2(new_n732), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n778), .A3(new_n785), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT110), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n994), .B1(new_n773), .B2(new_n992), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT109), .B1(new_n744), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1016), .A2(new_n996), .A3(new_n1029), .A4(new_n742), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n745), .B2(new_n996), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n744), .A2(new_n1027), .A3(KEYINPUT44), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n1008), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1023), .A2(new_n778), .A3(new_n785), .A4(KEYINPUT110), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1031), .A2(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(new_n740), .A3(new_n1034), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1026), .A2(new_n1040), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1012), .B1(new_n1044), .B2(new_n787), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n790), .B(KEYINPUT111), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1011), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n842), .A2(G68), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n818), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n882), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n260), .B1(new_n832), .B2(new_n349), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(KEYINPUT113), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(KEYINPUT113), .B2(new_n1052), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n829), .A2(new_n295), .B1(new_n880), .B2(new_n837), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT114), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n822), .A2(G143), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G50), .A2(new_n823), .B1(new_n820), .B2(G159), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT112), .B1(new_n830), .B2(G116), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT46), .Z(new_n1061));
  AOI21_X1  g0861(.A(new_n260), .B1(new_n834), .B2(G317), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n502), .B2(new_n826), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n832), .A2(new_n499), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G303), .C2(new_n818), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G283), .A2(new_n823), .B1(new_n822), .B2(G311), .ZN(new_n1066));
  INV_X1    g0866(.A(G294), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1066), .C1(new_n1067), .C2(new_n883), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1054), .A2(new_n1059), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT47), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n808), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n813), .B1(new_n747), .B2(new_n517), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n236), .A2(new_n800), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n793), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1073), .B(new_n1076), .C1(new_n857), .C2(new_n1004), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1048), .A2(new_n1077), .ZN(G387));
  AND2_X1   g0878(.A1(new_n1024), .A2(new_n748), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n787), .B2(new_n1023), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n800), .B1(new_n241), .B2(new_n491), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n751), .B2(new_n795), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n347), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n1083), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT50), .B1(new_n1083), .B2(G50), .ZN(new_n1085));
  AOI21_X1  g0885(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1084), .A2(new_n751), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1082), .A2(new_n1087), .B1(new_n502), .B2(new_n747), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n792), .B1(new_n1088), .B2(new_n813), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G50), .A2(new_n818), .B1(new_n822), .B2(G159), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n438), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G68), .A2(new_n823), .B1(new_n820), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n830), .A2(new_n222), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n826), .A2(new_n351), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n260), .B1(new_n837), .B2(new_n882), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1064), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n260), .B1(new_n834), .B2(G326), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n829), .A2(new_n1067), .B1(new_n826), .B2(new_n844), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G303), .A2(new_n823), .B1(new_n818), .B2(G317), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G311), .A2(new_n820), .B1(new_n822), .B2(G322), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT48), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1103), .B2(new_n1102), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT49), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1098), .B1(new_n647), .B2(new_n832), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1097), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1089), .B1(new_n1109), .B2(new_n808), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n737), .A2(new_n738), .A3(new_n811), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1023), .A2(new_n1047), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1080), .A2(new_n1112), .ZN(G393));
  NAND2_X1  g0913(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1024), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n1044), .A3(new_n748), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n996), .A2(new_n857), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT115), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n246), .A2(new_n801), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n813), .B1(G97), .B2(new_n747), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n820), .A2(G303), .B1(G116), .B2(new_n842), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT118), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n830), .A2(G283), .B1(G322), .B2(new_n834), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(KEYINPUT117), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(KEYINPUT117), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n258), .B1(new_n502), .B2(new_n832), .C1(new_n845), .C2(new_n1067), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G311), .A2(new_n818), .B1(new_n822), .B2(G317), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT52), .Z(new_n1130));
  AOI22_X1  g0930(.A1(G150), .A2(new_n822), .B1(new_n818), .B2(G159), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT51), .Z(new_n1132));
  OAI22_X1  g0932(.A1(new_n202), .A2(new_n883), .B1(new_n845), .B2(new_n1083), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT116), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n830), .A2(G68), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n842), .A2(G77), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n258), .B1(new_n834), .B2(G143), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n893), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1135), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1128), .A2(new_n1130), .B1(new_n1132), .B2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n792), .B1(new_n1119), .B2(new_n1121), .C1(new_n1142), .C2(new_n876), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1118), .A2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n1047), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1116), .A2(new_n1146), .ZN(G390));
  NAND3_X1  g0947(.A1(new_n716), .A2(new_n741), .A3(new_n869), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n867), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n869), .C1(new_n775), .C2(new_n777), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n953), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n731), .B1(new_n966), .B2(new_n970), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n954), .B1(new_n1153), .B2(new_n869), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n953), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n983), .A2(G330), .A3(new_n869), .A4(new_n954), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1150), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n698), .A2(new_n699), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n766), .A2(new_n967), .A3(KEYINPUT31), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n481), .B(G330), .C1(new_n775), .C2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1164), .A3(new_n959), .A4(new_n328), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT121), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n700), .A2(KEYINPUT121), .A3(new_n959), .A4(new_n1164), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1159), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT39), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n976), .A2(new_n922), .A3(new_n924), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT38), .B1(new_n1173), .B2(new_n911), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n943), .A2(new_n944), .A3(new_n927), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n945), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1176), .A2(new_n1177), .B1(new_n955), .B2(new_n948), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1175), .B1(new_n927), .B2(new_n926), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n953), .B1(new_n1148), .B2(new_n867), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n947), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT119), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n942), .A2(new_n946), .B1(new_n947), .B2(new_n1180), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n955), .A2(new_n948), .A3(new_n978), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1157), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1182), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1182), .A2(new_n1186), .A3(KEYINPUT120), .A4(new_n1187), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1183), .B(new_n1185), .C1(new_n953), .C2(new_n1151), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1171), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(new_n1192), .A3(new_n1191), .A4(new_n1170), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n748), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n809), .B1(new_n942), .B2(new_n946), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n792), .B1(new_n877), .B2(new_n1091), .ZN(new_n1199));
  INV_X1    g0999(.A(G125), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n260), .B1(new_n826), .B2(new_n838), .C1(new_n1200), .C2(new_n837), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n832), .A2(new_n202), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G137), .C2(new_n820), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT54), .B(G143), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n823), .A2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G128), .A2(new_n822), .B1(new_n818), .B2(G132), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n829), .A2(new_n882), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT53), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT122), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1138), .B(new_n258), .C1(new_n1067), .C2(new_n837), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G87), .B2(new_n830), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G107), .A2(new_n820), .B1(new_n818), .B2(G116), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G97), .A2(new_n823), .B1(new_n822), .B2(G283), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n887), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1210), .A2(KEYINPUT122), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1199), .B1(new_n1218), .B2(new_n808), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1198), .A2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n1047), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1197), .A2(new_n1222), .ZN(G378));
  XNOR2_X1  g1023(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n325), .A2(new_n918), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n329), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n329), .A2(new_n1227), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1225), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1225), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n809), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n792), .B1(new_n877), .B2(G50), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n818), .A2(G128), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n845), .B2(new_n880), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n830), .A2(new_n1205), .B1(G150), .B2(new_n842), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1200), .B2(new_n881), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G132), .C2(new_n820), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n833), .A2(G159), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n834), .C2(G124), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n502), .A2(new_n1050), .B1(new_n881), .B2(new_n647), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n499), .A2(new_n883), .B1(new_n845), .B2(new_n351), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n833), .A2(G58), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n258), .A2(new_n548), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G283), .B2(new_n834), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1093), .A2(new_n1250), .A3(new_n1049), .A4(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1248), .A2(new_n1249), .A3(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1251), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1247), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1236), .B1(new_n1258), .B2(new_n808), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1235), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1234), .B1(new_n981), .B2(new_n731), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1234), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n971), .A2(new_n980), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT40), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n971), .B2(new_n978), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G330), .B(new_n1262), .C1(new_n1264), .C2(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1261), .A2(new_n958), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n958), .B1(new_n1261), .B2(new_n1267), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1260), .B1(new_n1270), .B2(new_n1046), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1169), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1196), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1269), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1261), .A2(new_n958), .A3(new_n1267), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n748), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1270), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT57), .B1(new_n1274), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1272), .B1(new_n1280), .B2(new_n1282), .ZN(G375));
  OAI21_X1  g1083(.A(new_n792), .B1(new_n877), .B2(G68), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n260), .B(new_n1094), .C1(G303), .C2(new_n834), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1285), .B1(new_n345), .B2(new_n832), .C1(new_n499), .C2(new_n829), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(G283), .A2(new_n818), .B1(new_n822), .B2(G294), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1287), .B1(new_n502), .B2(new_n845), .C1(new_n647), .C2(new_n883), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(G132), .A2(new_n822), .B1(new_n818), .B2(G137), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n1289), .B1(new_n882), .B2(new_n845), .C1(new_n883), .C2(new_n1204), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n830), .A2(G159), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n842), .A2(G50), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n258), .B1(new_n834), .B2(G128), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1250), .A2(new_n1291), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n1286), .A2(new_n1288), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1284), .B1(new_n1295), .B2(new_n808), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n954), .B2(new_n810), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1159), .B2(new_n1046), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT123), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1012), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1159), .A2(new_n1169), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1171), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(G381));
  NOR3_X1   g1103(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1304), .A2(KEYINPUT124), .ZN(new_n1305));
  INV_X1    g1105(.A(G390), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(KEYINPUT124), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1308), .A2(G387), .A3(G381), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1197), .A2(new_n1222), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1274), .A2(new_n1281), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1275), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n749), .B1(new_n1274), .B2(new_n1278), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1271), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1309), .A2(new_n1310), .A3(new_n1314), .ZN(G407));
  INV_X1    g1115(.A(G213), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1316), .A2(G343), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1310), .A3(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(G407), .A2(G213), .A3(new_n1318), .ZN(G409));
  OAI211_X1 g1119(.A(G378), .B(new_n1272), .C1(new_n1280), .C2(new_n1282), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1272), .B1(new_n1311), .B2(new_n1012), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1310), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1317), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1301), .B1(new_n1170), .B2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1159), .A2(new_n1169), .A3(KEYINPUT60), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n748), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1299), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(G384), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1299), .A2(new_n1328), .A3(G384), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1323), .A2(new_n1324), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT62), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1317), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1338), .A2(new_n1339), .A3(new_n1334), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1317), .A2(G2897), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1331), .A2(new_n1332), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1341), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1270), .B1(new_n1196), .B2(new_n1273), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1271), .B1(new_n1346), .B2(new_n1300), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1347), .A2(G378), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1314), .B2(G378), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1345), .B1(new_n1349), .B2(new_n1317), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1336), .A2(new_n1337), .A3(new_n1340), .A4(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1044), .A2(new_n787), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1047), .B1(new_n1352), .B2(new_n1300), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1007), .B(new_n1009), .ZN(new_n1354));
  OAI211_X1 g1154(.A(G390), .B(new_n1077), .C1(new_n1353), .C2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT125), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(G387), .A2(new_n1306), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(G393), .A2(G396), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n859), .B1(new_n1080), .B2(new_n1112), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1048), .A2(KEYINPUT125), .A3(new_n1077), .A4(G390), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1357), .A2(new_n1358), .A3(new_n1362), .A4(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1364), .A2(KEYINPUT126), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1361), .B1(G387), .B2(new_n1306), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT126), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1366), .A2(new_n1367), .A3(new_n1357), .A4(new_n1363), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1365), .A2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1358), .A2(new_n1355), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1370), .A2(new_n1361), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1351), .A2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1341), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1333), .A2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1376), .A2(new_n1342), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1372), .B(new_n1337), .C1(new_n1338), .C2(new_n1377), .ZN(new_n1378));
  INV_X1    g1178(.A(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT63), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1335), .A2(new_n1380), .ZN(new_n1381));
  OAI21_X1  g1181(.A(KEYINPUT127), .B1(new_n1335), .B2(new_n1380), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT127), .ZN(new_n1383));
  NAND4_X1  g1183(.A1(new_n1338), .A2(new_n1383), .A3(KEYINPUT63), .A4(new_n1334), .ZN(new_n1384));
  NAND4_X1  g1184(.A1(new_n1379), .A2(new_n1381), .A3(new_n1382), .A4(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1374), .A2(new_n1385), .ZN(G405));
  NAND2_X1  g1186(.A1(G375), .A2(new_n1310), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1387), .A2(new_n1320), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1388), .A2(new_n1334), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1387), .A2(new_n1320), .A3(new_n1333), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1389), .A2(new_n1390), .ZN(new_n1391));
  XNOR2_X1  g1191(.A(new_n1391), .B(new_n1373), .ZN(G402));
endmodule


