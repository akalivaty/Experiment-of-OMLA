//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n190), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(G146), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT0), .A4(G128), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n189), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n201));
  OAI211_X1 g015(.A(G128), .B(new_n201), .C1(new_n193), .C2(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n197), .B(new_n198), .C1(KEYINPUT1), .C2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G125), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G224), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G953), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n200), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n207), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(new_n204), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n189), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n191), .A2(new_n190), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n199), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n208), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G116), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(G119), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n219), .A2(G119), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT2), .A2(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT2), .A3(G113), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT2), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n226), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n223), .A2(new_n231), .A3(new_n234), .A4(new_n225), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G104), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n239), .B2(G107), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  INV_X1    g055(.A(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(G107), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT76), .A2(G101), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT76), .A2(G101), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(new_n240), .A3(new_n243), .A4(new_n244), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(KEYINPUT4), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n252), .A3(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n238), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(G110), .B(G122), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n242), .A2(G104), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n244), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n256), .A2(new_n249), .B1(G101), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n223), .A2(KEYINPUT5), .A3(new_n225), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n233), .B1(new_n224), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n263), .A3(new_n237), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n254), .A2(new_n255), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n255), .A2(KEYINPUT81), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AND4_X1   g081(.A1(new_n234), .A2(new_n223), .A3(new_n231), .A4(new_n225), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n225), .A2(new_n223), .B1(new_n231), .B2(new_n234), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n253), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n251), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT80), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n254), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n276), .B2(KEYINPUT6), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n254), .A2(new_n274), .A3(new_n264), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n274), .B1(new_n254), .B2(new_n264), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT6), .B(new_n266), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n218), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n208), .B2(new_n216), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n200), .B2(new_n205), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n265), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n262), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n260), .B2(KEYINPUT82), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT69), .B(G116), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n224), .B1(new_n291), .B2(G119), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT82), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT5), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n237), .A3(new_n259), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n258), .A2(G101), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n237), .A2(new_n250), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n294), .B2(new_n290), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT83), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n228), .A2(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n260), .A2(new_n262), .B1(new_n292), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT84), .B1(new_n304), .B2(new_n259), .ZN(new_n305));
  INV_X1    g119(.A(new_n259), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n263), .A2(new_n237), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n298), .A2(new_n302), .A3(new_n305), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n255), .B(KEYINPUT8), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n288), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n283), .B1(new_n312), .B2(G902), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n305), .B(new_n309), .C1(new_n301), .C2(KEYINPUT83), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n296), .A2(new_n297), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n286), .A2(new_n265), .A3(new_n287), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G902), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(KEYINPUT85), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n282), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n322));
  OAI21_X1  g136(.A(G210), .B1(G237), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n321), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n282), .A2(new_n313), .A3(new_n323), .A4(new_n320), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT87), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n265), .A3(new_n280), .ZN(new_n333));
  AOI21_X1  g147(.A(G902), .B1(new_n316), .B2(new_n317), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n333), .A2(new_n218), .B1(new_n334), .B2(KEYINPUT85), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT87), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n323), .A4(new_n313), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n188), .B1(new_n327), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n203), .A2(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(KEYINPUT23), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT73), .B1(new_n340), .B2(G128), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G110), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n347), .A2(new_n352), .A3(KEYINPUT75), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n189), .A2(G140), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT16), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n189), .A2(G140), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT16), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(G146), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n358), .A2(G125), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n194), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n357), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n343), .A2(new_n344), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT72), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n361), .A2(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n194), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n365), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n350), .A2(new_n351), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G137), .ZN(new_n379));
  INV_X1    g193(.A(G953), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n380), .A2(G221), .A3(G234), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n379), .B(new_n381), .Z(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n369), .B1(new_n355), .B2(new_n356), .ZN(new_n385));
  INV_X1    g199(.A(new_n378), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(G234), .B2(new_n319), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n387), .A3(new_n319), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT25), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n383), .A2(new_n387), .A3(KEYINPUT25), .A4(new_n319), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n393), .B1(new_n398), .B2(new_n390), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(G472), .A2(G902), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n403));
  NOR2_X1   g217(.A1(G237), .A2(G953), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G210), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(G101), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n238), .ZN(new_n410));
  OR2_X1    g224(.A1(KEYINPUT64), .A2(G137), .ZN(new_n411));
  NAND2_X1  g225(.A1(KEYINPUT64), .A2(G137), .ZN(new_n412));
  AND2_X1   g226(.A1(KEYINPUT11), .A2(G134), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G137), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G134), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G134), .ZN(new_n419));
  AOI21_X1  g233(.A(G131), .B1(new_n419), .B2(G137), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n412), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(new_n419), .ZN(new_n424));
  INV_X1    g238(.A(G131), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(new_n210), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n419), .A2(G137), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n414), .A2(new_n418), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT65), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n429), .A2(new_n430), .A3(G131), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n429), .B2(G131), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n421), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n214), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n427), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n409), .B1(new_n410), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n414), .A2(new_n418), .A3(new_n420), .ZN(new_n438));
  AND2_X1   g252(.A1(KEYINPUT64), .A2(G137), .ZN(new_n439));
  NOR2_X1   g253(.A1(KEYINPUT64), .A2(G137), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n419), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n425), .B1(new_n441), .B2(new_n416), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n437), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n421), .B(KEYINPUT66), .C1(new_n424), .C2(new_n425), .ZN(new_n444));
  INV_X1    g258(.A(new_n210), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n434), .A2(new_n433), .B1(new_n446), .B2(KEYINPUT67), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT67), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n443), .A2(new_n448), .A3(new_n444), .A4(new_n445), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT30), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n433), .A2(new_n434), .ZN(new_n451));
  INV_X1    g265(.A(new_n427), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT30), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n238), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n436), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n451), .A2(new_n458), .A3(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n410), .B1(new_n435), .B2(KEYINPUT30), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT31), .A3(new_n436), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n410), .A3(new_n452), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT28), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT28), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n435), .A2(new_n468), .A3(new_n410), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n459), .A2(new_n238), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n409), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n402), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n463), .A2(new_n475), .A3(new_n466), .A4(new_n409), .ZN(new_n476));
  INV_X1    g290(.A(new_n469), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n468), .B1(new_n435), .B2(new_n410), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n471), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n408), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n435), .A2(new_n410), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n475), .B1(new_n470), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n319), .B(new_n476), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n474), .A2(KEYINPUT32), .B1(G472), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n408), .B1(new_n470), .B2(new_n471), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n457), .B2(new_n464), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n487), .B2(new_n402), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n400), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n367), .B(new_n194), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n380), .A3(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n192), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n404), .A2(G143), .A3(G214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT18), .A3(G131), .ZN(new_n496));
  AND4_X1   g310(.A1(G143), .A2(new_n491), .A3(new_n380), .A4(G214), .ZN(new_n497));
  AOI21_X1  g311(.A(G143), .B1(new_n404), .B2(G214), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n425), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n497), .B2(new_n498), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n495), .A2(KEYINPUT88), .A3(G131), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n499), .A2(new_n425), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n361), .A2(G146), .A3(new_n364), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n362), .B2(new_n366), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n511), .ZN(new_n514));
  NAND2_X1  g328(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n359), .A3(new_n360), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G146), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n510), .B1(new_n517), .B2(KEYINPUT90), .ZN(new_n518));
  AND4_X1   g332(.A1(new_n359), .A2(new_n514), .A3(new_n360), .A4(new_n515), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT19), .B1(new_n359), .B2(new_n360), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n194), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n509), .B1(new_n524), .B2(KEYINPUT91), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n518), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n503), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n239), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT92), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(G146), .B1(new_n361), .B2(new_n364), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT93), .B1(new_n510), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n375), .A2(new_n534), .A3(new_n365), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT88), .B1(new_n495), .B2(G131), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n505), .B(new_n425), .C1(new_n493), .C2(new_n494), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT17), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n536), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n530), .A3(new_n502), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n542), .A2(KEYINPUT94), .A3(new_n530), .A4(new_n502), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n512), .A2(new_n516), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT90), .A3(new_n194), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n365), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n517), .A2(KEYINPUT90), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT91), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n509), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n527), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n502), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n556));
  INV_X1    g370(.A(new_n530), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n531), .A2(new_n547), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT20), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n531), .A2(new_n547), .A3(new_n558), .A4(KEYINPUT95), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n562), .B1(new_n566), .B2(KEYINPUT20), .ZN(new_n567));
  INV_X1    g381(.A(G475), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n542), .A2(new_n502), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n557), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n547), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n571), .B2(new_n319), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT9), .B(G234), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n573), .A2(new_n389), .A3(G953), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT13), .B1(new_n203), .B2(G143), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n419), .ZN(new_n576));
  XNOR2_X1  g390(.A(G128), .B(G143), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n291), .A2(G122), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n219), .A2(G122), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n242), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n242), .B1(new_n579), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n577), .B(new_n419), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT14), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n579), .A2(new_n586), .A3(new_n580), .ZN(new_n587));
  OAI21_X1  g401(.A(G107), .B1(new_n579), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n581), .B(new_n585), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n574), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n584), .A2(new_n589), .A3(new_n574), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n593), .A2(new_n319), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n591), .B2(new_n592), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n600), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n319), .B(new_n380), .C1(G234), .C2(G237), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT21), .B(G898), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n380), .A2(G952), .ZN(new_n609));
  INV_X1    g423(.A(G234), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n491), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n567), .A2(new_n572), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n573), .B2(G902), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n251), .A2(new_n434), .A3(new_n253), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n250), .A2(new_n204), .A3(new_n202), .A4(new_n299), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n619), .A2(KEYINPUT77), .A3(KEYINPUT10), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT10), .B1(new_n619), .B2(KEYINPUT77), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT78), .B1(new_n622), .B2(new_n433), .ZN(new_n623));
  INV_X1    g437(.A(new_n621), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n619), .A2(KEYINPUT77), .A3(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT78), .ZN(new_n627));
  INV_X1    g441(.A(new_n433), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n618), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n306), .A2(new_n210), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n619), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n433), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT12), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(KEYINPUT12), .A3(new_n433), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(G110), .B(G140), .ZN(new_n639));
  INV_X1    g453(.A(G227), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(G953), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n623), .B2(new_n629), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n626), .A2(KEYINPUT79), .A3(new_n618), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT79), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n646), .A3(new_n433), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n638), .A2(new_n642), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(G469), .B1(new_n648), .B2(G902), .ZN(new_n649));
  INV_X1    g463(.A(G469), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n643), .A2(new_n637), .ZN(new_n651));
  INV_X1    g465(.A(new_n642), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n630), .B2(new_n647), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n650), .B(new_n319), .C1(new_n651), .C2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n617), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n339), .A2(new_n489), .A3(new_n615), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(new_n249), .Z(G3));
  NAND2_X1  g472(.A1(new_n603), .A2(new_n594), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n594), .A2(new_n319), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT99), .B1(new_n593), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n663), .A2(KEYINPUT33), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT33), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n593), .B2(KEYINPUT99), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n659), .B(new_n661), .C1(new_n668), .C2(new_n594), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n566), .A2(KEYINPUT20), .ZN(new_n670));
  INV_X1    g484(.A(new_n562), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n545), .A2(new_n546), .B1(new_n557), .B2(new_n569), .ZN(new_n673));
  OAI21_X1  g487(.A(G475), .B1(new_n673), .B2(G902), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n669), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n321), .A2(new_n324), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n612), .B(new_n188), .C1(new_n676), .C2(new_n328), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(KEYINPUT100), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n659), .A2(new_n661), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n664), .A2(new_n667), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(G478), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n567), .B2(new_n572), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n188), .B1(new_n676), .B2(new_n328), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n613), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n679), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n649), .A2(new_n654), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n399), .A3(new_n616), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n487), .B2(G902), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n463), .A2(KEYINPUT31), .A3(new_n436), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT31), .B1(new_n463), .B2(new_n436), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n473), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n401), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT34), .B(G104), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G6));
  NOR2_X1   g513(.A1(new_n572), .A2(new_n605), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n613), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n564), .A2(new_n560), .A3(new_n561), .A4(new_n565), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n670), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n684), .B1(new_n703), .B2(KEYINPUT101), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n705), .B(new_n701), .C1(new_n670), .C2(new_n702), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n696), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT35), .B(G107), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G9));
  NAND2_X1  g524(.A1(new_n371), .A2(new_n378), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n384), .A2(KEYINPUT36), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n711), .B(new_n712), .Z(new_n713));
  AOI22_X1  g527(.A1(new_n398), .A2(new_n390), .B1(new_n713), .B2(new_n391), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n695), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n339), .A2(new_n615), .A3(new_n655), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT37), .B(G110), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G12));
  NAND2_X1  g532(.A1(new_n483), .A2(G472), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n693), .A2(KEYINPUT32), .A3(new_n401), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n488), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n714), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n655), .A3(new_n684), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n606), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n611), .B1(new_n724), .B2(G900), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT102), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n670), .B2(new_n702), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n700), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n203), .ZN(G30));
  NAND2_X1  g544(.A1(new_n676), .A2(KEYINPUT86), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n338), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT38), .Z(new_n734));
  XOR2_X1   g548(.A(new_n726), .B(KEYINPUT39), .Z(new_n735));
  NAND2_X1  g549(.A1(new_n655), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT40), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n722), .A2(new_n605), .A3(new_n188), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n672), .A2(new_n674), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n481), .A2(new_n466), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n409), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT103), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n741), .A2(KEYINPUT103), .B1(new_n463), .B2(new_n436), .ZN(new_n743));
  AOI21_X1  g557(.A(G902), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(G472), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n488), .B(new_n720), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n738), .A2(new_n739), .A3(new_n746), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n734), .A2(new_n737), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  INV_X1    g563(.A(new_n726), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n682), .B(new_n750), .C1(new_n567), .C2(new_n572), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n714), .B1(new_n484), .B2(new_n488), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n684), .A2(new_n655), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT104), .B1(new_n723), .B2(new_n751), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G146), .ZN(G48));
  NAND2_X1  g573(.A1(new_n630), .A2(new_n647), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n760), .A2(new_n642), .B1(new_n643), .B2(new_n637), .ZN(new_n761));
  OAI21_X1  g575(.A(G469), .B1(new_n761), .B2(G902), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n616), .A3(new_n654), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n721), .A2(new_n399), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n678), .B2(new_n686), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT41), .B(G113), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G15));
  NOR3_X1   g582(.A1(new_n704), .A2(new_n706), .A3(new_n765), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n219), .ZN(G18));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n567), .A2(new_n572), .ZN(new_n772));
  INV_X1    g586(.A(new_n614), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n684), .A4(new_n764), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n721), .A2(new_n722), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n676), .A2(new_n328), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n187), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n763), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n753), .A2(new_n779), .A3(KEYINPUT105), .A4(new_n615), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G119), .ZN(G21));
  NOR2_X1   g596(.A1(new_n763), .A2(new_n612), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n470), .A2(new_n481), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n465), .B1(new_n408), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n401), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n783), .A2(new_n399), .A3(new_n690), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n605), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n684), .B(new_n788), .C1(new_n572), .C2(new_n567), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(G122), .Z(G24));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n739), .A2(new_n792), .A3(new_n682), .A4(new_n750), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n786), .A2(new_n690), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n714), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n779), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G125), .ZN(G27));
  NAND4_X1  g612(.A1(new_n338), .A2(new_n731), .A3(new_n187), .A4(new_n732), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT107), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n648), .B2(G469), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n617), .B1(new_n803), .B2(new_n654), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT32), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n694), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n400), .B1(new_n484), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n793), .A2(new_n806), .A3(new_n794), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n751), .B(new_n792), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n327), .A2(new_n187), .A3(new_n338), .A4(new_n804), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n721), .A2(new_n399), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(KEYINPUT42), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g628(.A1(KEYINPUT42), .A2(new_n810), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G131), .ZN(G33));
  NOR3_X1   g630(.A1(new_n812), .A2(new_n813), .A3(new_n728), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n419), .ZN(G36));
  NOR2_X1   g632(.A1(new_n648), .A2(KEYINPUT45), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n650), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n648), .A2(KEYINPUT45), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n801), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT46), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n654), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n799), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n616), .A3(new_n735), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n772), .A2(new_n682), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT43), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT108), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT43), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n831), .B(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT108), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n714), .B1(new_n690), .B2(new_n694), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT44), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n830), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT44), .A4(new_n838), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G137), .ZN(G39));
  OR4_X1    g658(.A1(new_n721), .A2(new_n751), .A3(new_n799), .A4(new_n399), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n828), .A2(KEYINPUT47), .A3(new_n616), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n616), .B1(new_n826), .B2(new_n827), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n358), .ZN(G42));
  OR4_X1    g665(.A1(new_n400), .A2(new_n831), .A3(new_n617), .A4(new_n188), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT109), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n762), .A2(new_n654), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT49), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n746), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n853), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n857), .A3(new_n734), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n339), .A2(new_n613), .A3(new_n696), .A4(new_n675), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n656), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n567), .A2(new_n572), .A3(new_n605), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n733), .A3(new_n613), .A4(new_n187), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n339), .A2(KEYINPUT111), .A3(new_n613), .A4(new_n864), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n696), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n869), .A3(new_n716), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n766), .A2(new_n769), .A3(new_n790), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT110), .B1(new_n872), .B2(new_n781), .ZN(new_n873));
  INV_X1    g687(.A(new_n765), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n790), .B1(new_n707), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n687), .A2(new_n874), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n781), .A4(KEYINPUT110), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n871), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n729), .ZN(new_n880));
  INV_X1    g694(.A(new_n789), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n805), .A2(new_n722), .A3(new_n726), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n746), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n758), .A2(new_n880), .A3(new_n797), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT52), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n793), .A2(new_n794), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n829), .A2(new_n809), .A3(new_n804), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT42), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n812), .A2(new_n813), .ZN(new_n889));
  INV_X1    g703(.A(new_n728), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n674), .A2(new_n605), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n617), .B(new_n891), .C1(new_n649), .C2(new_n654), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n721), .A2(new_n727), .A3(new_n892), .A4(new_n722), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n889), .A2(new_n890), .B1(new_n893), .B2(new_n829), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n811), .A2(new_n814), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n888), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT112), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n829), .A2(new_n796), .A3(new_n804), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n886), .B2(new_n898), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n799), .A2(new_n795), .A3(new_n805), .A4(new_n714), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(KEYINPUT112), .A3(new_n794), .A4(new_n793), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n729), .B1(new_n756), .B2(new_n757), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n797), .A4(new_n883), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n885), .A2(new_n896), .A3(new_n902), .A4(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n861), .B1(new_n879), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n875), .A2(new_n876), .A3(new_n781), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT110), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n870), .B1(new_n910), .B2(new_n877), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n885), .A2(new_n905), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n902), .A2(new_n815), .A3(new_n894), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT53), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n860), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n867), .A2(new_n868), .A3(new_n696), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n656), .A2(new_n716), .A3(new_n862), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n861), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n875), .A2(new_n876), .A3(new_n781), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n896), .A4(new_n902), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n885), .A2(new_n905), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT113), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT113), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n863), .A2(new_n869), .A3(KEYINPUT53), .A4(new_n716), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n908), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n912), .A2(new_n924), .A3(new_n914), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n923), .A2(new_n927), .B1(new_n928), .B2(new_n861), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n916), .B1(new_n860), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n832), .A2(new_n611), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n795), .A2(new_n400), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n763), .A2(new_n187), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT114), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n734), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT50), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n846), .B(new_n849), .C1(new_n616), .C2(new_n855), .ZN(new_n939));
  INV_X1    g753(.A(new_n933), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n829), .A3(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n746), .A2(new_n400), .A3(new_n611), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n799), .A2(new_n763), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n944), .A2(new_n739), .A3(new_n682), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n931), .A2(new_n943), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n796), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n938), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n940), .A2(new_n779), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n609), .C1(new_n683), .C2(new_n944), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n946), .A2(new_n809), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT48), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT115), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(KEYINPUT115), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n953), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AND4_X1   g774(.A1(new_n930), .A2(new_n950), .A3(new_n951), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(G952), .A2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n859), .B1(new_n961), .B2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n380), .A2(G952), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n913), .A2(new_n908), .A3(new_n925), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n924), .B1(new_n965), .B2(new_n912), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n921), .A2(KEYINPUT113), .A3(new_n922), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n907), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(G210), .A3(G902), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT56), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n333), .B(new_n217), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT55), .Z(new_n973));
  AOI21_X1  g787(.A(new_n964), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT116), .ZN(new_n975));
  INV_X1    g789(.A(new_n973), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n969), .A2(new_n975), .A3(new_n970), .A4(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n969), .A2(new_n970), .A3(new_n976), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(KEYINPUT116), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(G51));
  XOR2_X1   g794(.A(new_n801), .B(KEYINPUT57), .Z(new_n981));
  NOR2_X1   g795(.A1(new_n968), .A2(KEYINPUT54), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n923), .A2(new_n927), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n860), .B1(new_n983), .B2(new_n907), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n653), .B2(new_n651), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n822), .B(KEYINPUT117), .Z(new_n987));
  NAND3_X1  g801(.A1(new_n968), .A2(G902), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n964), .B1(new_n986), .B2(new_n988), .ZN(G54));
  INV_X1    g803(.A(KEYINPUT118), .ZN(new_n990));
  INV_X1    g804(.A(new_n964), .ZN(new_n991));
  NAND2_X1  g805(.A1(KEYINPUT58), .A2(G475), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n319), .B(new_n992), .C1(new_n983), .C2(new_n907), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n564), .A2(new_n565), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n968), .A2(G902), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n997), .A2(new_n994), .A3(new_n992), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n990), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n993), .A2(new_n995), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n994), .B1(new_n997), .B2(new_n992), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT118), .A4(new_n991), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(G60));
  XNOR2_X1  g817(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n661), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n681), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n982), .B2(new_n984), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n991), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n929), .A2(new_n860), .ZN(new_n1010));
  INV_X1    g824(.A(new_n916), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT120), .B1(new_n1012), .B2(new_n668), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT120), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1014), .B(new_n681), .C1(new_n930), .C2(new_n1006), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1009), .B1(new_n1013), .B2(new_n1015), .ZN(G63));
  XNOR2_X1  g830(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(G217), .A2(G902), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT60), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n968), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n388), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n991), .ZN(new_n1024));
  INV_X1    g838(.A(new_n713), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1018), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n964), .B1(new_n1022), .B2(new_n388), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1028), .B(new_n1017), .C1(new_n1025), .C2(new_n1022), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(G66));
  OAI21_X1  g844(.A(G953), .B1(new_n607), .B2(new_n206), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n911), .B2(G953), .ZN(new_n1032));
  INV_X1    g846(.A(new_n333), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(G898), .B2(new_n380), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT124), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1032), .B(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g850(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(G69));
  AOI21_X1  g852(.A(new_n850), .B1(new_n841), .B2(new_n842), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n903), .A2(new_n797), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n748), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT62), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1040), .A2(KEYINPUT62), .A3(new_n748), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n813), .A2(new_n799), .A3(new_n736), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1046), .B1(new_n675), .B2(new_n864), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1039), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n380), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n461), .A2(new_n453), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1050), .B(new_n548), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n881), .A2(new_n809), .ZN(new_n1053));
  INV_X1    g867(.A(new_n735), .ZN(new_n1054));
  NOR3_X1   g868(.A1(new_n847), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n1055), .A2(new_n817), .ZN(new_n1056));
  AND3_X1   g870(.A1(new_n1056), .A2(new_n1040), .A3(new_n815), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1039), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(KEYINPUT125), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1039), .A2(KEYINPUT125), .A3(new_n1057), .ZN(new_n1061));
  AND3_X1   g875(.A1(new_n1060), .A2(new_n380), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1051), .ZN(new_n1063));
  INV_X1    g877(.A(G900), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1063), .B1(new_n1064), .B2(new_n380), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1052), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g880(.A(G953), .B1(new_n640), .B2(new_n1064), .C1(new_n1051), .C2(KEYINPUT126), .ZN(new_n1067));
  INV_X1    g881(.A(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g882(.A(new_n1066), .B(new_n1068), .ZN(G72));
  INV_X1    g883(.A(KEYINPUT127), .ZN(new_n1070));
  NAND2_X1  g884(.A1(G472), .A2(G902), .ZN(new_n1071));
  XOR2_X1   g885(.A(new_n1071), .B(KEYINPUT63), .Z(new_n1072));
  OAI21_X1  g886(.A(new_n1072), .B1(new_n1048), .B2(new_n879), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n409), .B1(new_n463), .B2(new_n466), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n964), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n907), .A2(new_n915), .ZN(new_n1076));
  NAND3_X1  g890(.A1(new_n463), .A2(new_n466), .A3(new_n409), .ZN(new_n1077));
  INV_X1    g891(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g892(.A(new_n1072), .ZN(new_n1079));
  NOR3_X1   g893(.A1(new_n1078), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1080));
  NAND2_X1  g894(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g895(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g896(.A1(new_n1060), .A2(new_n911), .A3(new_n1061), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n1077), .B1(new_n1083), .B2(new_n1072), .ZN(new_n1084));
  OAI21_X1  g898(.A(new_n1070), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1083), .A2(new_n1072), .ZN(new_n1086));
  NAND2_X1  g900(.A1(new_n1086), .A2(new_n1078), .ZN(new_n1087));
  NAND4_X1  g901(.A1(new_n1087), .A2(KEYINPUT127), .A3(new_n1081), .A4(new_n1075), .ZN(new_n1088));
  NAND2_X1  g902(.A1(new_n1085), .A2(new_n1088), .ZN(G57));
endmodule


