//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT68), .A3(G119), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G116), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n190), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n192), .A3(G116), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT68), .B1(new_n187), .B2(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(new_n189), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT69), .B1(new_n201), .B2(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(G104), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n204), .A2(new_n211), .A3(new_n205), .A4(G104), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n208), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT5), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT86), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT86), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT5), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n219), .B1(new_n224), .B2(new_n189), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n201), .B2(new_n224), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n203), .A2(new_n218), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n207), .A2(new_n210), .A3(new_n212), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n231), .A3(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n198), .A2(new_n202), .B1(new_n201), .B2(new_n196), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n227), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT87), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n227), .B(new_n236), .C1(new_n233), .C2(new_n234), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n235), .A2(KEYINPUT6), .A3(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT0), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT65), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(KEYINPUT0), .B2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n249), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(G125), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n255), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n256), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n254), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n254), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n260), .A2(new_n255), .A3(new_n257), .A4(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n262), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n259), .B(KEYINPUT88), .C1(G125), .C2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(KEYINPUT88), .B2(new_n259), .ZN(new_n272));
  INV_X1    g086(.A(G224), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G953), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n272), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n243), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n195), .B1(new_n194), .B2(new_n197), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n201), .A2(KEYINPUT69), .A3(new_n196), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n217), .B(new_n226), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n236), .B(KEYINPUT8), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT5), .B(new_n199), .C1(new_n200), .C2(new_n189), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n198), .A2(new_n202), .B1(new_n225), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n280), .B(new_n281), .C1(new_n217), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n275), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n259), .B(KEYINPUT90), .C1(G125), .C2(new_n270), .ZN(new_n288));
  OR3_X1    g102(.A1(new_n270), .A2(KEYINPUT90), .A3(G125), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n275), .A2(KEYINPUT7), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT91), .A4(new_n290), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n286), .A2(new_n287), .A3(new_n295), .A4(new_n241), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n277), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n243), .B2(new_n276), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n299), .A3(new_n296), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT84), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT85), .Z(new_n307));
  NAND2_X1  g121(.A1(G234), .A2(G237), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(G952), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT21), .B(G898), .Z(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(G902), .A3(G953), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n307), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT9), .B(G234), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G221), .B1(new_n320), .B2(G902), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT78), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G469), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(G137), .ZN(new_n329));
  INV_X1    g143(.A(G137), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT11), .A3(G134), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n331), .A3(new_n334), .A4(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n262), .A2(new_n269), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n217), .A3(new_n267), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n270), .A2(new_n213), .A3(new_n216), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n325), .B1(new_n341), .B2(KEYINPUT12), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT12), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n217), .B(new_n270), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT82), .B(new_n343), .C1(new_n344), .C2(new_n337), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n348));
  INV_X1    g162(.A(new_n251), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n258), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n230), .A2(new_n350), .A3(new_n232), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n218), .A2(KEYINPUT10), .A3(new_n270), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n351), .A2(new_n353), .A3(new_n354), .A4(new_n337), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n309), .A2(G227), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT79), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G140), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(KEYINPUT80), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(KEYINPUT80), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n347), .A2(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n361), .A2(new_n355), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n336), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT83), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n347), .A2(new_n355), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n368), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n324), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n347), .A2(new_n365), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(new_n355), .ZN(new_n378));
  INV_X1    g192(.A(new_n361), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n324), .A3(new_n297), .ZN(new_n382));
  NAND2_X1  g196(.A1(G469), .A2(G902), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n323), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n318), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n330), .A2(G134), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n327), .A2(G137), .ZN(new_n388));
  OAI21_X1  g202(.A(G131), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n335), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n336), .A2(new_n350), .B1(new_n270), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT67), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n350), .A2(new_n336), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n270), .A2(new_n390), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT67), .ZN(new_n397));
  INV_X1    g211(.A(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI22_X1  g213(.A1(new_n278), .A2(new_n279), .B1(new_n194), .B2(new_n197), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(KEYINPUT30), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n393), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT70), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT26), .B(G101), .Z(new_n405));
  NOR2_X1   g219(.A1(G237), .A2(G953), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G210), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n405), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n391), .A2(new_n234), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n404), .A2(KEYINPUT31), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n413));
  AOI211_X1 g227(.A(KEYINPUT67), .B(new_n392), .C1(new_n394), .C2(new_n395), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n403), .A3(new_n400), .A4(new_n401), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n410), .A3(new_n411), .A4(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n396), .A2(new_n400), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n391), .A2(new_n234), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT28), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT28), .B1(new_n391), .B2(new_n234), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n410), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT31), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G472), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n412), .A2(new_n427), .A3(new_n428), .A4(new_n297), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n418), .B2(new_n426), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT32), .A3(new_n412), .A4(new_n428), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n421), .A2(KEYINPUT29), .A3(new_n410), .A4(new_n423), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n396), .A2(new_n400), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n411), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n422), .B1(new_n438), .B2(KEYINPUT28), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n439), .A2(KEYINPUT72), .A3(KEYINPUT29), .A4(new_n410), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n416), .A2(new_n411), .A3(new_n417), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n442), .B2(new_n425), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n410), .ZN(new_n444));
  AOI211_X1 g258(.A(G902), .B(new_n441), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n431), .B(new_n433), .C1(new_n445), .C2(new_n428), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT22), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(G137), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT76), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n360), .A3(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n360), .A2(G125), .ZN(new_n453));
  INV_X1    g267(.A(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(G146), .B(new_n452), .C1(new_n456), .C2(new_n451), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT74), .ZN(new_n458));
  XNOR2_X1  g272(.A(G125), .B(G140), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT16), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT74), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G146), .A4(new_n452), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n192), .B2(G128), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n192), .A2(G128), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n245), .A2(KEYINPUT23), .A3(G119), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n358), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n245), .A2(G119), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n466), .B2(new_n470), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT24), .B(G110), .Z(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n459), .A2(new_n254), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n463), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n479));
  INV_X1    g293(.A(new_n477), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n458), .B2(new_n462), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n476), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n468), .A2(new_n358), .ZN(new_n485));
  INV_X1    g299(.A(new_n472), .ZN(new_n486));
  INV_X1    g300(.A(new_n473), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n475), .ZN(new_n488));
  INV_X1    g302(.A(new_n457), .ZN(new_n489));
  AOI21_X1  g303(.A(G146), .B1(new_n460), .B2(new_n452), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n450), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  AOI211_X1 g307(.A(KEYINPUT76), .B(new_n493), .C1(new_n479), .C2(new_n483), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n449), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n479), .B2(new_n483), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n449), .B1(new_n496), .B2(new_n450), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT77), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n495), .A2(new_n297), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n499), .A2(KEYINPUT77), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND4_X1   g317(.A1(new_n482), .A2(new_n463), .A3(new_n476), .A4(new_n477), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n482), .B1(new_n481), .B2(new_n476), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n491), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT76), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n484), .A2(new_n450), .A3(new_n491), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n497), .B1(new_n509), .B2(new_n449), .ZN(new_n510));
  INV_X1    g324(.A(new_n502), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n510), .A2(new_n297), .A3(new_n511), .A4(new_n500), .ZN(new_n512));
  INV_X1    g326(.A(G217), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(G234), .B2(new_n297), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(G902), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G475), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n406), .A2(G143), .A3(G214), .ZN(new_n521));
  AOI21_X1  g335(.A(G143), .B1(new_n406), .B2(G214), .ZN(new_n522));
  OAI21_X1  g336(.A(G131), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT93), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n525), .B(G131), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT97), .B1(new_n489), .B2(new_n490), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n521), .A2(new_n522), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n334), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n524), .A2(new_n531), .A3(new_n532), .A4(new_n526), .ZN(new_n533));
  INV_X1    g347(.A(new_n490), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n457), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n528), .A2(new_n529), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n456), .A2(G146), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n477), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n530), .B1(KEYINPUT18), .B2(G131), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n530), .A2(KEYINPUT18), .A3(G131), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(G113), .B(G122), .Z(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT96), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(new_n214), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n537), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n537), .B2(new_n544), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n520), .B1(new_n550), .B2(new_n297), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n524), .A2(new_n526), .A3(new_n531), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n553));
  OR3_X1    g367(.A1(new_n456), .A2(new_n553), .A3(KEYINPUT95), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT95), .B1(new_n456), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n456), .A2(KEYINPUT19), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n552), .B(new_n463), .C1(G146), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n544), .ZN(new_n559));
  INV_X1    g373(.A(new_n547), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n537), .A2(new_n544), .A3(new_n547), .ZN(new_n562));
  AOI21_X1  g376(.A(G475), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n297), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n563), .B2(new_n297), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(KEYINPUT98), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n562), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n520), .A3(new_n297), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n569), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n551), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n245), .A2(G143), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n263), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n327), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n245), .B2(G143), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n263), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(KEYINPUT13), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(new_n579), .C1(new_n577), .C2(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G134), .ZN(new_n581));
  XNOR2_X1  g395(.A(G116), .B(G122), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT99), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n205), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(new_n205), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n574), .B(new_n581), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(KEYINPUT101), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n573), .B(new_n327), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n583), .A2(new_n590), .A3(new_n205), .ZN(new_n591));
  INV_X1    g405(.A(G122), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(new_n592), .B2(G116), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n187), .B2(G122), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n592), .A2(KEYINPUT14), .A3(G116), .ZN(new_n595));
  OAI21_X1  g409(.A(G107), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n319), .A2(G217), .A3(new_n309), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n587), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G478), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n603), .A2(new_n606), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n571), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n386), .A2(new_n446), .A3(new_n519), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  NAND2_X1  g428(.A1(new_n432), .A2(new_n412), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G472), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n429), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n518), .ZN(new_n618));
  INV_X1    g432(.A(new_n385), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT102), .ZN(new_n621));
  INV_X1    g435(.A(new_n551), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT98), .B1(new_n569), .B2(KEYINPUT20), .ZN(new_n623));
  INV_X1    g437(.A(new_n565), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n569), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n600), .A2(new_n602), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n600), .A2(KEYINPUT33), .A3(new_n602), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n630), .A2(G478), .A3(new_n297), .A4(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n603), .A2(G478), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n306), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n297), .A2(new_n277), .A3(new_n299), .A4(new_n296), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n299), .B1(new_n302), .B2(new_n296), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n637), .B(new_n317), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n621), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT34), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n214), .ZN(G6));
  INV_X1    g458(.A(new_n609), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n607), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n646), .B(new_n622), .C1(new_n624), .C2(new_n566), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n621), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT104), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT35), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G107), .ZN(G9));
  INV_X1    g465(.A(new_n617), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n506), .B(KEYINPUT105), .ZN(new_n653));
  INV_X1    g467(.A(new_n449), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n516), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n515), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n386), .A2(new_n612), .A3(new_n652), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AND2_X1   g475(.A1(new_n431), .A2(new_n433), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n443), .A2(new_n444), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n297), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n664), .B2(new_n441), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n385), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n306), .B1(new_n301), .B2(new_n303), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n658), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n311), .B1(new_n315), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n647), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n666), .A2(KEYINPUT106), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n446), .A2(new_n619), .A3(new_n672), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n675), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n671), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n619), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n658), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n304), .B(KEYINPUT38), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n571), .A2(new_n610), .A3(new_n306), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n425), .B1(new_n404), .B2(new_n411), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n297), .B1(new_n438), .B2(new_n410), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n662), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n682), .A2(new_n685), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NAND2_X1  g506(.A1(new_n567), .A2(new_n570), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n634), .B1(new_n693), .B2(new_n622), .ZN(new_n694));
  INV_X1    g508(.A(new_n671), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n571), .A2(new_n634), .A3(new_n671), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT107), .B1(new_n700), .B2(new_n667), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n658), .B(new_n666), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NOR2_X1   g517(.A1(new_n636), .A2(new_n640), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n347), .A2(new_n365), .B1(new_n378), .B2(new_n379), .ZN(new_n705));
  OAI21_X1  g519(.A(G469), .B1(new_n705), .B2(G902), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n382), .A3(new_n323), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n704), .A2(new_n446), .A3(new_n519), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT108), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n709), .B(new_n711), .ZN(G15));
  NOR2_X1   g526(.A1(new_n640), .A2(new_n647), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n446), .A2(new_n713), .A3(new_n519), .A4(new_n708), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n698), .B2(new_n707), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n667), .A2(KEYINPUT109), .A3(new_n708), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n611), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n446), .A3(new_n317), .A4(new_n658), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  AOI21_X1  g535(.A(new_n316), .B1(new_n301), .B2(new_n303), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n618), .A2(new_n722), .A3(new_n684), .A4(new_n708), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n515), .A2(new_n657), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n725), .B1(new_n726), .B2(new_n617), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n658), .A2(KEYINPUT110), .A3(new_n429), .A4(new_n616), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n696), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n717), .A2(new_n718), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND3_X1  g546(.A1(new_n373), .A2(G469), .A3(new_n368), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n382), .A2(new_n733), .A3(new_n383), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n323), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n301), .A2(new_n637), .A3(new_n303), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n446), .A2(new_n519), .A3(new_n700), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT42), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n334), .ZN(G33));
  INV_X1    g554(.A(new_n446), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n518), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n672), .A3(new_n737), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  NAND3_X1  g558(.A1(new_n373), .A2(KEYINPUT45), .A3(new_n368), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n370), .A2(new_n375), .ZN(new_n746));
  OAI211_X1 g560(.A(G469), .B(new_n745), .C1(new_n746), .C2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n383), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n383), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n382), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n323), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n679), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT111), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(KEYINPUT111), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n635), .A2(new_n571), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n652), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n758), .B(KEYINPUT43), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n726), .B1(new_n763), .B2(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n736), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT113), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n762), .A2(new_n764), .A3(new_n769), .A4(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n757), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n753), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n753), .A2(new_n775), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n753), .A2(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n753), .A2(new_n775), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n696), .A2(new_n519), .A3(new_n736), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n741), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  AND2_X1   g599(.A1(new_n706), .A2(new_n382), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n322), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n778), .A2(new_n781), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n736), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n760), .A2(new_n311), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(KEYINPUT121), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n760), .B2(new_n311), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n618), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n788), .A2(new_n789), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n519), .A2(new_n311), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n789), .A2(new_n708), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n689), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n571), .A3(new_n634), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT123), .Z(new_n802));
  OAI21_X1  g616(.A(KEYINPUT122), .B1(new_n794), .B2(new_n799), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n790), .B(KEYINPUT121), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n805));
  INV_X1    g619(.A(new_n799), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n727), .A2(new_n728), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n802), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n618), .A3(new_n708), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n683), .A2(new_n637), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n796), .A2(KEYINPUT50), .A3(new_n708), .A4(new_n813), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n797), .A2(new_n810), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(G952), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n821), .B(G953), .C1(new_n800), .C2(new_n694), .ZN(new_n822));
  INV_X1    g636(.A(new_n742), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n803), .B2(new_n807), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n822), .B1(new_n824), .B2(KEYINPUT48), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(KEYINPUT48), .B2(new_n824), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n797), .A2(new_n810), .A3(new_n817), .A4(KEYINPUT51), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n796), .A2(new_n730), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n684), .A2(new_n304), .ZN(new_n830));
  INV_X1    g644(.A(new_n735), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n671), .B(KEYINPUT119), .Z(new_n832));
  NOR2_X1   g646(.A1(new_n658), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n689), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n677), .A2(KEYINPUT118), .A3(new_n731), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT118), .B1(new_n677), .B2(new_n731), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n702), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n720), .A2(new_n709), .A3(new_n714), .A4(new_n723), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n739), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT115), .B1(new_n636), .B2(new_n318), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n694), .A2(new_n843), .A3(new_n307), .A4(new_n722), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n619), .A3(new_n618), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n610), .A2(KEYINPUT116), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n646), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n627), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n386), .A2(new_n618), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n845), .A2(new_n613), .A3(new_n659), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n737), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n696), .B(new_n853), .C1(new_n727), .C2(new_n728), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n624), .A2(new_n566), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n551), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n849), .A2(new_n856), .A3(new_n695), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n789), .B1(new_n857), .B2(KEYINPUT117), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n849), .A2(new_n856), .A3(KEYINPUT117), .A4(new_n695), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n446), .A3(new_n619), .A4(new_n658), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n852), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n677), .A2(new_n702), .A3(new_n731), .A4(new_n834), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n862), .B(new_n743), .C1(new_n863), .C2(KEYINPUT52), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n841), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT53), .B1(new_n868), .B2(new_n864), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n840), .B2(new_n739), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n738), .B(new_n874), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n446), .A2(new_n713), .A3(new_n519), .A4(new_n708), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n611), .B(new_n726), .C1(new_n718), .C2(new_n717), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n741), .A2(new_n316), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n709), .A2(new_n723), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT120), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n882), .B(new_n864), .C1(KEYINPUT52), .C2(new_n837), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n839), .B1(new_n868), .B2(new_n864), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n828), .A2(new_n829), .A3(new_n871), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n821), .A2(new_n309), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n683), .A2(new_n518), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n635), .A2(new_n571), .A3(new_n323), .A4(new_n307), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n786), .B(KEYINPUT49), .Z(new_n894));
  OR4_X1    g708(.A1(new_n689), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(G75));
  XNOR2_X1  g710(.A(KEYINPUT124), .B(KEYINPUT55), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n243), .B(new_n276), .Z(new_n898));
  INV_X1    g712(.A(new_n882), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n838), .A2(new_n865), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n297), .B1(new_n900), .B2(new_n884), .ZN(new_n901));
  AOI211_X1 g715(.A(KEYINPUT56), .B(new_n898), .C1(new_n901), .C2(G210), .ZN(new_n902));
  INV_X1    g716(.A(new_n898), .ZN(new_n903));
  OAI211_X1 g717(.A(G210), .B(G902), .C1(new_n883), .C2(new_n885), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n309), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(G210), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n910), .B(new_n297), .C1(new_n900), .C2(new_n884), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n898), .B1(new_n911), .B2(KEYINPUT56), .ZN(new_n912));
  INV_X1    g726(.A(new_n897), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n904), .A2(new_n905), .A3(new_n903), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n907), .A2(new_n909), .A3(new_n915), .ZN(G51));
  NAND2_X1  g730(.A1(new_n900), .A2(new_n884), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n887), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n383), .B(KEYINPUT57), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n381), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n886), .A2(new_n297), .A3(new_n747), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND3_X1  g736(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n923));
  INV_X1    g737(.A(new_n568), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n908), .ZN(G60));
  NAND2_X1  g741(.A1(new_n630), .A2(new_n631), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n871), .A2(new_n888), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n932), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n935), .A3(new_n908), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n886), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n656), .ZN(new_n940));
  INV_X1    g754(.A(new_n510), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n886), .B2(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n909), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n909), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(G66));
  OR2_X1    g761(.A1(new_n840), .A2(new_n852), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n309), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n313), .B2(new_n273), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n243), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(G898), .B2(new_n309), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G69));
  INV_X1    g768(.A(G227), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n955), .B2(new_n670), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n784), .A2(new_n875), .A3(new_n743), .A4(new_n772), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n835), .A2(new_n836), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n702), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n757), .A2(new_n742), .A3(new_n830), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n309), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n670), .A2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n415), .A2(new_n401), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n557), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n959), .A2(new_n691), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n446), .B1(new_n778), .B2(new_n781), .ZN(new_n969));
  AOI22_X1  g783(.A1(new_n755), .A2(new_n756), .B1(new_n768), .B2(new_n770), .ZN(new_n970));
  AOI22_X1  g784(.A1(new_n969), .A2(new_n783), .B1(new_n970), .B2(new_n767), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n958), .A2(new_n691), .A3(new_n702), .ZN(new_n972));
  XNOR2_X1  g786(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n680), .A2(new_n736), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n975), .B(new_n742), .C1(new_n694), .C2(new_n850), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n968), .A2(new_n971), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n965), .A2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(KEYINPUT127), .B(new_n956), .C1(new_n966), .C2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n982));
  AND4_X1   g796(.A1(new_n981), .A2(new_n966), .A3(new_n982), .A4(new_n979), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n980), .A2(new_n983), .ZN(G72));
  NOR2_X1   g798(.A1(new_n442), .A2(new_n410), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n957), .A2(new_n961), .A3(new_n948), .ZN(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n686), .A2(new_n985), .A3(new_n989), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n870), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n909), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n988), .B1(new_n977), .B2(new_n948), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n686), .B2(new_n994), .ZN(G57));
endmodule


