//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G131), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G134), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G137), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT11), .B1(new_n190), .B2(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G134), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(KEYINPUT67), .A3(new_n189), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n192), .B2(G137), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(new_n198), .A3(new_n189), .A4(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n194), .B1(new_n199), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(G146), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(G146), .B1(new_n212), .B2(new_n214), .ZN(new_n219));
  AOI21_X1  g033(.A(G143), .B1(new_n207), .B2(new_n209), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n216), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n205), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n201), .A2(new_n198), .A3(new_n193), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n199), .A2(new_n204), .B1(G131), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n219), .B2(new_n220), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n210), .A2(new_n215), .A3(KEYINPUT0), .A4(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT2), .B(G113), .Z(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n225), .A2(G131), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n202), .A2(new_n203), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n202), .A2(new_n203), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n231), .A2(new_n232), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n205), .A2(new_n223), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(new_n238), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n242), .B(new_n252), .C1(new_n239), .C2(new_n235), .ZN(new_n253));
  INV_X1    g067(.A(G237), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G210), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT27), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n259), .B(KEYINPUT69), .Z(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n259), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT30), .B1(new_n224), .B2(new_n234), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n248), .A2(new_n265), .A3(new_n249), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT68), .B1(new_n267), .B2(new_n238), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n269), .B(new_n239), .C1(new_n264), .C2(new_n266), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n240), .B(new_n263), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n262), .B1(new_n271), .B2(KEYINPUT31), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n248), .A2(new_n265), .A3(new_n249), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n265), .B1(new_n248), .B2(new_n249), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n238), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n269), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n267), .A2(KEYINPUT68), .A3(new_n238), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n251), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n273), .B1(new_n279), .B2(new_n263), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n187), .B(new_n188), .C1(new_n272), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n271), .A2(KEYINPUT31), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n273), .A3(new_n263), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n262), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n188), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n253), .B2(new_n261), .ZN(new_n289));
  INV_X1    g103(.A(new_n279), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n259), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT71), .B1(new_n235), .B2(new_n239), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n250), .A2(new_n293), .A3(new_n238), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n251), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n242), .B1(new_n295), .B2(new_n241), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n188), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G472), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n283), .A2(new_n287), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT79), .ZN(new_n302));
  OAI21_X1  g116(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n246), .A2(KEYINPUT80), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n226), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT10), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n210), .A2(new_n215), .A3(new_n217), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n210), .A2(new_n215), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n312));
  OAI21_X1  g126(.A(G128), .B1(new_n219), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G104), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(new_n315), .B2(G107), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G104), .ZN(new_n319));
  INV_X1    g133(.A(G101), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(G107), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n316), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n315), .A2(G107), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n318), .A2(G104), .ZN(new_n324));
  OAI21_X1  g138(.A(G101), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n309), .B1(new_n314), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n319), .A3(new_n321), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G101), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n331), .A3(G101), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n232), .A3(new_n231), .A4(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n326), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n308), .A2(new_n327), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n226), .A2(KEYINPUT81), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n313), .A2(new_n311), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n326), .B1(new_n338), .B2(new_n218), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n218), .B(new_n326), .C1(new_n221), .C2(new_n222), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n340), .B1(new_n314), .B2(new_n326), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT12), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n337), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G140), .ZN(new_n348));
  INV_X1    g162(.A(G227), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n348), .B(new_n350), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n335), .B(new_n333), .C1(new_n339), .C2(KEYINPUT10), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n246), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n336), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT82), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(G469), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G469), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n336), .A2(new_n343), .A3(new_n351), .A4(new_n346), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n351), .B1(new_n355), .B2(new_n336), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n362), .B(new_n188), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(G469), .A2(G902), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n304), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G478), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT15), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n302), .A2(new_n371), .A3(G953), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G116), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(G116), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n212), .A2(new_n214), .A3(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n216), .A2(G143), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n192), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n318), .B1(new_n376), .B2(new_n377), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT90), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT65), .B(G143), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(KEYINPUT91), .A3(KEYINPUT13), .A4(G128), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n380), .A2(new_n390), .A3(new_n385), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n381), .A2(KEYINPUT91), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n380), .B2(new_n385), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n387), .A2(new_n389), .A3(new_n391), .A4(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n394), .B2(G134), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n318), .B1(new_n375), .B2(KEYINPUT14), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n378), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n380), .A2(new_n381), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G134), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n382), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n373), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n400), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n380), .A2(new_n385), .ZN(new_n404));
  AOI22_X1  g218(.A1(KEYINPUT91), .A2(new_n404), .B1(new_n386), .B2(KEYINPUT90), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT13), .B1(new_n388), .B2(G128), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(KEYINPUT13), .A3(G128), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n406), .A2(new_n390), .B1(new_n407), .B2(new_n392), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n192), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n403), .B(new_n372), .C1(new_n409), .C2(new_n384), .ZN(new_n410));
  AOI21_X1  g224(.A(G902), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n370), .B1(new_n411), .B2(KEYINPUT92), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n188), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(KEYINPUT92), .A3(new_n370), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G140), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G125), .ZN(new_n421));
  INV_X1    g235(.A(G125), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G140), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT16), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n422), .A2(KEYINPUT16), .A3(G140), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n206), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n425), .A3(new_n428), .A4(G146), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n254), .A2(new_n255), .A3(G214), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n212), .A3(new_n214), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n254), .A2(new_n255), .A3(G143), .A4(G214), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n189), .A3(new_n433), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n424), .A2(new_n425), .A3(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n189), .B1(new_n432), .B2(new_n433), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n430), .A2(new_n438), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(new_n315), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT66), .B(G146), .ZN(new_n446));
  XNOR2_X1  g260(.A(G125), .B(G140), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n206), .B2(new_n447), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n189), .ZN(new_n451));
  OAI221_X1 g265(.A(new_n449), .B1(new_n434), .B2(new_n451), .C1(new_n435), .C2(new_n450), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n443), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n445), .B1(new_n443), .B2(new_n452), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n188), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n454), .B(new_n445), .C1(new_n443), .C2(new_n452), .ZN(new_n458));
  OAI21_X1  g272(.A(G475), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n432), .A2(new_n189), .A3(new_n433), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT87), .B1(new_n460), .B2(new_n441), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n435), .A2(new_n462), .A3(new_n437), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n421), .A2(new_n423), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n447), .A2(KEYINPUT19), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n422), .A2(KEYINPUT16), .A3(G140), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n468), .A2(new_n446), .B1(G146), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT88), .A3(new_n452), .ZN(new_n473));
  INV_X1    g287(.A(new_n445), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT88), .B1(new_n472), .B2(new_n452), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n453), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n459), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G952), .ZN(new_n483));
  AOI211_X1 g297(.A(G953), .B(new_n483), .C1(G234), .C2(G237), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n188), .B(new_n255), .C1(G234), .C2(G237), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(G898), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n419), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G214), .B1(G237), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT85), .B1(new_n326), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n237), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g307(.A(G116), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(KEYINPUT5), .A3(G119), .ZN(new_n495));
  INV_X1    g309(.A(G113), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n493), .A2(new_n497), .B1(new_n236), .B2(new_n237), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n492), .B(new_n499), .C1(KEYINPUT85), .C2(new_n326), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n498), .B(KEYINPUT85), .C1(new_n491), .C2(new_n326), .ZN(new_n501));
  XNOR2_X1  g315(.A(G110), .B(G122), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT8), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n238), .A2(new_n330), .A3(new_n332), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n334), .A2(new_n498), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n223), .A2(new_n422), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n231), .A2(G125), .A3(new_n232), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n255), .A2(G224), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT7), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n504), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n312), .B1(new_n446), .B2(G143), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n515), .A2(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n516));
  AOI21_X1  g330(.A(G125), .B1(new_n516), .B2(new_n218), .ZN(new_n517));
  INV_X1    g331(.A(new_n509), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(KEYINPUT86), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n505), .A2(new_n506), .ZN(new_n525));
  INV_X1    g339(.A(new_n502), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT83), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n507), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n508), .A2(new_n510), .A3(new_n509), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n510), .B1(new_n508), .B2(new_n509), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n525), .B(new_n526), .C1(KEYINPUT83), .C2(new_n528), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G210), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n524), .A2(new_n537), .A3(new_n535), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n490), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n368), .A2(new_n488), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n371), .B1(G234), .B2(new_n188), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT75), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n440), .A2(new_n429), .A3(new_n427), .ZN(new_n545));
  XOR2_X1   g359(.A(G119), .B(G128), .Z(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT24), .B(G110), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT23), .B1(new_n216), .B2(G119), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n216), .A2(G119), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n216), .B(G119), .C1(KEYINPUT72), .C2(KEYINPUT23), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n548), .B1(new_n554), .B2(G110), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n546), .A2(new_n547), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n554), .B2(G110), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n439), .A2(new_n448), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND4_X1   g377(.A1(new_n544), .A2(new_n556), .A3(new_n559), .A4(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n545), .A2(new_n555), .B1(new_n561), .B2(new_n562), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n544), .B1(new_n565), .B2(new_n559), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n556), .A2(new_n563), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT74), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n559), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n567), .A2(KEYINPUT25), .A3(new_n573), .A4(new_n188), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n567), .A2(new_n188), .A3(new_n573), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n577));
  AOI22_X1  g391(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n575), .A3(new_n577), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n543), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n543), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n567), .A2(new_n188), .A3(new_n573), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT78), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n300), .A2(new_n542), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AND2_X1   g400(.A1(new_n584), .A2(new_n368), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n281), .A2(KEYINPUT93), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n187), .B1(new_n286), .B2(new_n188), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(KEYINPUT93), .B(new_n187), .C1(new_n286), .C2(new_n188), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT94), .B(new_n587), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n524), .A2(new_n537), .A3(new_n535), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n537), .B1(new_n524), .B2(new_n535), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n489), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n599), .A2(new_n487), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n410), .A2(KEYINPUT95), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n413), .A2(new_n601), .A3(KEYINPUT33), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n402), .B(new_n410), .C1(KEYINPUT95), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n369), .A2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n414), .A2(KEYINPUT96), .A3(new_n369), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n411), .B2(G478), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n482), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n600), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n596), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NAND2_X1  g432(.A1(new_n417), .A2(new_n418), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n600), .A2(new_n482), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n596), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT98), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NAND2_X1  g438(.A1(new_n569), .A2(new_n571), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n188), .A3(new_n581), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n580), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n368), .A2(new_n488), .A3(new_n629), .A4(new_n541), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n590), .B2(new_n591), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G12));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n484), .B1(new_n485), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n482), .A2(new_n619), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n368), .A2(new_n541), .A3(new_n629), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n300), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  XOR2_X1   g453(.A(new_n635), .B(KEYINPUT39), .Z(new_n640));
  NAND2_X1  g454(.A1(new_n368), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n539), .A2(new_n540), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n419), .A2(new_n482), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n489), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n647), .A3(new_n629), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n271), .B1(new_n260), .B2(new_n295), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n188), .B1(new_n649), .B2(new_n650), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n287), .A3(new_n283), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n642), .A2(new_n648), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(new_n388), .Z(G45));
  INV_X1    g471(.A(new_n635), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n482), .A2(new_n612), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n368), .A2(new_n660), .A3(new_n629), .A4(new_n541), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n300), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT101), .B(G146), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G48));
  OAI21_X1  g478(.A(new_n188), .B1(new_n363), .B2(new_n364), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G469), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n303), .A3(new_n365), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n300), .A2(new_n668), .A3(new_n584), .A4(new_n614), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  NAND4_X1  g485(.A1(new_n300), .A2(new_n620), .A3(new_n584), .A4(new_n668), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G116), .ZN(G18));
  NOR2_X1   g487(.A1(new_n667), .A2(new_n599), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n488), .A3(new_n629), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n300), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G119), .ZN(G21));
  NOR2_X1   g491(.A1(new_n667), .A2(new_n487), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n541), .A2(new_n482), .A3(new_n419), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(KEYINPUT103), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n646), .B2(new_n541), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n188), .B1(new_n272), .B2(new_n280), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n296), .A2(new_n261), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n284), .A2(new_n285), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(G472), .A2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n584), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n584), .A4(new_n689), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n683), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n374), .ZN(G24));
  INV_X1    g509(.A(new_n688), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n251), .B(new_n259), .C1(new_n277), .C2(new_n278), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n697), .A2(new_n273), .B1(new_n261), .B2(new_n296), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n698), .B2(new_n284), .ZN(new_n699));
  INV_X1    g513(.A(new_n628), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n576), .A2(new_n575), .A3(new_n577), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n574), .A2(new_n575), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n576), .A2(new_n577), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(new_n704), .B2(new_n543), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n589), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n659), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n482), .A2(new_n612), .A3(KEYINPUT104), .A4(new_n658), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n709), .A2(new_n674), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n685), .A2(new_n629), .A3(new_n689), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(new_n674), .A3(new_n710), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  INV_X1    g531(.A(KEYINPUT32), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n281), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n287), .A3(new_n299), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n584), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n539), .A2(new_n303), .A3(new_n489), .A4(new_n540), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n365), .B(new_n366), .C1(new_n357), .C2(new_n362), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n709), .A2(new_n710), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT42), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n300), .A2(new_n584), .A3(new_n728), .A4(new_n727), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n721), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n189), .ZN(G33));
  NAND4_X1  g547(.A1(new_n300), .A2(new_n584), .A3(new_n636), .A4(new_n727), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  INV_X1    g549(.A(new_n612), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n482), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT108), .B1(new_n737), .B2(KEYINPUT43), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n738), .A2(new_n740), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n590), .A2(new_n591), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n629), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n539), .A2(new_n489), .A3(new_n540), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n747), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n358), .A2(new_n360), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n753));
  INV_X1    g567(.A(new_n357), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n362), .B1(new_n754), .B2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n366), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n365), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT46), .B1(new_n756), .B2(new_n366), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n303), .B(new_n640), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  OR4_X1    g577(.A1(new_n300), .A2(new_n584), .A3(new_n659), .A4(new_n749), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n303), .B1(new_n758), .B2(new_n759), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT47), .B(new_n303), .C1(new_n758), .C2(new_n759), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n420), .ZN(G42));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n666), .A2(new_n365), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n645), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n737), .A2(new_n303), .A3(new_n489), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(KEYINPUT49), .B2(new_n772), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n584), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n774), .B1(new_n777), .B2(KEYINPUT109), .ZN(new_n778));
  INV_X1    g592(.A(new_n654), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n778), .B(new_n779), .C1(KEYINPUT109), .C2(new_n777), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n744), .A2(new_n484), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n692), .A2(new_n693), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n674), .A3(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(G952), .A3(new_n255), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n722), .A2(new_n772), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n584), .A3(new_n484), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT117), .ZN(new_n787));
  INV_X1    g601(.A(new_n613), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n785), .ZN(new_n791));
  INV_X1    g605(.A(new_n721), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n784), .B(new_n789), .C1(new_n793), .C2(KEYINPUT48), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n781), .A2(KEYINPUT118), .A3(new_n721), .A4(new_n785), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT48), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n791), .A2(new_n713), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(KEYINPUT50), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n645), .A2(new_n490), .A3(new_n668), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT115), .Z(new_n803));
  NAND3_X1  g617(.A1(new_n781), .A2(new_n803), .A3(new_n782), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n798), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n482), .A2(new_n612), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n787), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n772), .B(KEYINPUT114), .Z(new_n808));
  OAI211_X1 g622(.A(new_n767), .B(new_n768), .C1(new_n303), .C2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n809), .A2(new_n750), .B1(new_n803), .B2(new_n800), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n781), .A2(new_n782), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n805), .B(new_n807), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n797), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n631), .A2(new_n585), .A3(new_n676), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n694), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n619), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n482), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n788), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n600), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n594), .A2(new_n595), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n672), .A2(new_n669), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n749), .A2(new_n482), .A3(new_n635), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n368), .A2(new_n826), .A3(new_n819), .A4(new_n629), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(KEYINPUT111), .A3(new_n300), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT111), .B1(new_n827), .B2(new_n300), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n721), .A2(new_n729), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n730), .A2(new_n731), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n706), .A2(new_n728), .A3(new_n727), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(new_n734), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n830), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n679), .B(KEYINPUT103), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n580), .A2(new_n303), .A3(new_n628), .A4(new_n658), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n726), .B2(new_n725), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n654), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n300), .B1(new_n661), .B2(new_n637), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n707), .B1(new_n706), .B2(new_n711), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT105), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n716), .A2(KEYINPUT52), .A3(new_n841), .A4(new_n842), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT53), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n851), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n817), .A2(new_n823), .A3(new_n824), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n734), .B(new_n834), .C1(new_n828), .C2(new_n829), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n732), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n837), .A2(new_n860), .A3(KEYINPUT53), .A4(new_n849), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n850), .A2(new_n852), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  MUX2_X1   g679(.A(new_n854), .B(new_n864), .S(new_n865), .Z(new_n866));
  AND2_X1   g680(.A1(new_n815), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n771), .B(new_n780), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n815), .B2(new_n866), .ZN(new_n870));
  INV_X1    g684(.A(new_n780), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(G75));
  NOR2_X1   g687(.A1(new_n255), .A2(G952), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n188), .B1(new_n862), .B2(new_n863), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT56), .B1(new_n876), .B2(G210), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n530), .A2(new_n534), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(new_n533), .Z(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n875), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n877), .B2(new_n880), .ZN(G51));
  NOR2_X1   g696(.A1(new_n363), .A2(new_n364), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n862), .A2(new_n865), .A3(new_n863), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n366), .B(KEYINPUT57), .Z(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n756), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n864), .A2(G902), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT120), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n876), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n875), .B1(new_n888), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(KEYINPUT121), .B(new_n875), .C1(new_n888), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(G54));
  AND2_X1   g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n876), .A2(new_n477), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n876), .A2(new_n900), .ZN(new_n905));
  INV_X1    g719(.A(new_n477), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n874), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT123), .A4(new_n904), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(G60));
  INV_X1    g726(.A(new_n605), .ZN(new_n913));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT59), .Z(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n866), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n874), .B1(new_n886), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(G63));
  OAI21_X1  g733(.A(KEYINPUT60), .B1(new_n371), .B2(new_n188), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n371), .A2(new_n188), .A3(KEYINPUT60), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n864), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n627), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n875), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT61), .B1(new_n924), .B2(KEYINPUT124), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n567), .A2(new_n573), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n927), .B(new_n875), .C1(new_n923), .C2(new_n922), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n925), .B(new_n928), .ZN(G66));
  NAND2_X1  g743(.A1(G224), .A2(G953), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n825), .A2(G953), .B1(new_n486), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(G898), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n878), .B1(new_n932), .B2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  XOR2_X1   g748(.A(new_n267), .B(new_n468), .Z(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT125), .Z(new_n936));
  AND2_X1   g750(.A1(new_n716), .A2(new_n842), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n656), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  INV_X1    g753(.A(new_n769), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n821), .A2(new_n641), .A3(new_n749), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n300), .A3(new_n584), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n939), .A2(new_n762), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n943), .B2(new_n255), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n255), .A2(G900), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n761), .A2(new_n838), .A3(new_n721), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n940), .A2(new_n734), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(new_n833), .A3(new_n762), .A4(new_n937), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n945), .B1(new_n948), .B2(new_n255), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n935), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n349), .B2(new_n634), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n943), .B2(new_n825), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n290), .A3(new_n263), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n279), .A2(new_n263), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n957), .B1(new_n960), .B2(new_n697), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n854), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n948), .A2(new_n825), .ZN(new_n963));
  INV_X1    g777(.A(new_n957), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n279), .A2(new_n259), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n875), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(G57));
endmodule


