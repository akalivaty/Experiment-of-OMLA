//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n207), .A2(new_n208), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n212), .ZN(new_n214));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n222), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n217), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G141gat), .B(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(G155gat), .B2(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n213), .A2(new_n216), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n229), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(KEYINPUT5), .A3(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n213), .A2(new_n216), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n236), .A2(new_n237), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n236), .A2(new_n237), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n236), .B2(new_n237), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT73), .B1(new_n252), .B2(new_n217), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT3), .B1(new_n227), .B2(new_n228), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n249), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n254), .A2(KEYINPUT73), .A3(new_n217), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n240), .B(new_n248), .C1(new_n253), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n247), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n217), .A3(new_n255), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(new_n256), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n259), .B1(new_n266), .B2(new_n240), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n242), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G57gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(KEYINPUT75), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT75), .ZN(new_n274));
  INV_X1    g073(.A(new_n242), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n240), .A3(new_n259), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n272), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n279), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n273), .A2(new_n280), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT6), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G8gat), .B(G36gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G64gat), .ZN(new_n288));
  INV_X1    g087(.A(G92gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G211gat), .A2(G218gat), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(KEYINPUT22), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(new_n291), .A3(new_n294), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n296), .A2(new_n297), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G226gat), .ZN(new_n305));
  INV_X1    g104(.A(G233gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n312), .A2(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT66), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G190gat), .ZN(new_n323));
  AOI21_X1  g122(.A(G183gat), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n314), .B(KEYINPUT25), .C1(new_n319), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT66), .B(G190gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(G183gat), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(KEYINPUT67), .A3(KEYINPUT25), .A4(new_n314), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT64), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n320), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n335), .B1(new_n340), .B2(new_n319), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n330), .A2(KEYINPUT65), .A3(new_n339), .A4(new_n338), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n314), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n310), .A2(new_n311), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(KEYINPUT26), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(KEYINPUT26), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n315), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT69), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G183gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT28), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n352), .B1(new_n356), .B2(new_n331), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n321), .A2(new_n323), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT69), .A4(KEYINPUT28), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OR3_X1    g161(.A1(new_n337), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT27), .B1(new_n337), .B2(KEYINPUT68), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n334), .A2(new_n345), .B1(new_n351), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n308), .B1(new_n369), .B2(KEYINPUT29), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n327), .A3(new_n333), .ZN(new_n371));
  INV_X1    g170(.A(new_n367), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n351), .B1(new_n372), .B2(new_n361), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n308), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n304), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n343), .A2(new_n344), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n327), .A2(new_n333), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n307), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n303), .B1(new_n301), .B2(KEYINPUT72), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n298), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n381), .A2(new_n383), .A3(new_n374), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n290), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n304), .A3(new_n375), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n381), .B2(new_n374), .ZN(new_n387));
  INV_X1    g186(.A(new_n290), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(KEYINPUT30), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(new_n387), .A3(new_n391), .A4(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n286), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n383), .B1(KEYINPUT29), .B2(new_n250), .ZN(new_n395));
  INV_X1    g194(.A(G228gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n306), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n304), .B2(new_n380), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n395), .B(new_n397), .C1(new_n398), .C2(new_n244), .ZN(new_n399));
  INV_X1    g198(.A(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n380), .B1(new_n382), .B2(new_n298), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n244), .B1(new_n401), .B2(new_n249), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n250), .A2(KEYINPUT29), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n304), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G22gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n399), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT31), .B(G50gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT76), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G78gat), .ZN(new_n413));
  INV_X1    g212(.A(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n407), .A2(new_n408), .A3(new_n410), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n415), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n399), .A2(new_n405), .A3(new_n409), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n409), .B1(new_n399), .B2(new_n405), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n416), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n394), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G71gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G99gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n371), .A2(new_n243), .A3(new_n373), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n243), .B1(new_n371), .B2(new_n373), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n379), .A2(new_n217), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n428), .B1(new_n436), .B2(new_n430), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT70), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n440), .A3(KEYINPUT32), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n433), .B(KEYINPUT32), .C1(new_n434), .C2(new_n427), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n436), .A2(new_n430), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(new_n429), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n436), .A2(KEYINPUT34), .A3(new_n428), .A4(new_n430), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n442), .A2(new_n450), .A3(new_n443), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT36), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(KEYINPUT71), .A3(new_n448), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n442), .A2(new_n443), .A3(new_n453), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT36), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n424), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n248), .B1(new_n253), .B2(new_n257), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT78), .A3(new_n241), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n266), .B2(new_n240), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n229), .A2(new_n240), .A3(new_n238), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n467), .A2(KEYINPUT39), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n466), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n462), .A2(new_n464), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT40), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT79), .B(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT78), .B1(new_n461), .B2(new_n241), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n266), .A2(new_n463), .A3(new_n240), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n272), .ZN(new_n479));
  INV_X1    g278(.A(new_n474), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n462), .B2(new_n464), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT80), .B1(new_n481), .B2(new_n279), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n473), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n392), .B(new_n390), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n486), .B(new_n473), .C1(new_n479), .C2(new_n482), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n485), .A2(new_n284), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT37), .B1(new_n376), .B2(new_n384), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n386), .A2(new_n387), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n290), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n389), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n489), .A2(new_n493), .A3(new_n290), .A4(new_n491), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(new_n283), .A3(new_n285), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n422), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n460), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n497), .A2(new_n422), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n479), .A2(new_n482), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n486), .B1(new_n501), .B2(new_n473), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n484), .ZN(new_n503));
  INV_X1    g302(.A(new_n393), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n282), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT83), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n459), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n422), .A2(new_n455), .A3(new_n456), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT84), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  AOI221_X4 g310(.A(new_n511), .B1(new_n390), .B2(new_n392), .C1(new_n283), .C2(new_n285), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n422), .A2(new_n455), .A3(KEYINPUT84), .A4(new_n456), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n286), .A2(new_n422), .A3(new_n393), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n449), .A2(new_n451), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n202), .B1(new_n507), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n459), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n500), .A2(KEYINPUT83), .A3(new_n505), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT83), .B1(new_n500), .B2(new_n505), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT85), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G183gat), .B(G211gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G1gat), .B2(new_n530), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G71gat), .B(G78gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G127gat), .B(G155gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n529), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  INV_X1    g351(.A(new_n529), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n541), .A2(new_n542), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n551), .A2(new_n554), .A3(new_n558), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT91), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT41), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT92), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G190gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G218gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT93), .B(G85gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n574), .A2(new_n289), .B1(KEYINPUT8), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT94), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G99gat), .B(G106gat), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n581), .A3(new_n579), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G29gat), .ZN(new_n586));
  INV_X1    g385(.A(G36gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT14), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT14), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(G29gat), .B2(G36gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n591), .A2(KEYINPUT86), .B1(G29gat), .B2(G36gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(KEYINPUT86), .B2(new_n591), .ZN(new_n593));
  XOR2_X1   g392(.A(G43gat), .B(G50gat), .Z(new_n594));
  INV_X1    g393(.A(KEYINPUT15), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT88), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(KEYINPUT87), .A3(new_n596), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n591), .B1(new_n595), .B2(new_n594), .ZN(new_n603));
  OAI221_X1 g402(.A(new_n603), .B1(new_n595), .B2(new_n594), .C1(new_n586), .C2(new_n587), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n604), .A2(KEYINPUT88), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT17), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n608), .A3(new_n605), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n585), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n599), .A2(new_n601), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n604), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n585), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n565), .B2(new_n564), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n573), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n610), .A2(new_n614), .A3(new_n573), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n570), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n569), .A3(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n562), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n602), .A2(new_n608), .A3(new_n605), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n608), .B1(new_n602), .B2(new_n605), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n535), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n535), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT18), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n611), .A2(new_n535), .A3(new_n604), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(KEYINPUT89), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n626), .B(KEYINPUT13), .Z(new_n634));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n612), .A2(new_n635), .A3(new_n627), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n625), .A2(KEYINPUT18), .A3(new_n626), .A4(new_n628), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT11), .B(G169gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G197gat), .ZN(new_n641));
  XOR2_X1   g440(.A(G113gat), .B(G141gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n631), .A2(new_n644), .A3(new_n637), .A4(new_n638), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n583), .A2(new_n541), .A3(new_n584), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n576), .A2(KEYINPUT94), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n576), .A2(KEYINPUT94), .ZN(new_n652));
  OAI211_X1 g451(.A(KEYINPUT97), .B(new_n579), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT98), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT97), .B1(new_n581), .B2(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n654), .A2(new_n581), .B1(new_n580), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n649), .B(new_n650), .C1(new_n657), .C2(new_n541), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n540), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n657), .A2(new_n541), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n650), .ZN(new_n664));
  INV_X1    g463(.A(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n311), .ZN(new_n668));
  INV_X1    g467(.A(G204gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n662), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n665), .B1(new_n658), .B2(new_n659), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n661), .B1(new_n663), .B2(new_n650), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT99), .B(new_n670), .C1(new_n673), .C2(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n648), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n622), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n526), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n286), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT100), .B(G1gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1324gat));
  NOR2_X1   g484(.A1(new_n682), .A2(new_n393), .ZN(new_n686));
  NAND2_X1  g485(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n531), .A2(new_n534), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n691), .B(new_n692), .C1(new_n534), .C2(new_n686), .ZN(G1325gat));
  INV_X1    g492(.A(new_n682), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n458), .A2(new_n452), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n694), .A2(G15gat), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n516), .ZN(new_n697));
  AOI21_X1  g496(.A(G15gat), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n422), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(new_n621), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n680), .A2(new_n562), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n519), .A2(new_n525), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n286), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n519), .A2(new_n525), .A3(new_n703), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n518), .A2(KEYINPUT103), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n514), .A2(new_n712), .A3(new_n517), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT44), .B1(new_n714), .B2(new_n523), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n619), .A2(new_n569), .A3(new_n615), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n569), .B1(new_n619), .B2(new_n615), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n618), .A2(new_n620), .A3(KEYINPUT104), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n710), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n704), .B(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n286), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n726), .ZN(G1328gat));
  OAI21_X1  g526(.A(G36gat), .B1(new_n725), .B2(new_n393), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n705), .A2(G36gat), .A3(new_n393), .ZN(new_n729));
  AND2_X1   g528(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n728), .B(new_n732), .C1(new_n730), .C2(new_n729), .ZN(G1329gat));
  NOR3_X1   g532(.A1(new_n705), .A2(G43gat), .A3(new_n516), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n723), .A2(new_n695), .A3(new_n724), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g537(.A(KEYINPUT47), .B(new_n734), .C1(new_n735), .C2(G43gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1330gat));
  NOR3_X1   g539(.A1(new_n705), .A2(G50gat), .A3(new_n422), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n423), .A3(new_n724), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(G50gat), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT48), .B(new_n741), .C1(new_n742), .C2(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1331gat));
  NAND2_X1  g546(.A1(new_n714), .A2(new_n523), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n622), .A2(new_n648), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n677), .A2(new_n678), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n286), .B(KEYINPUT106), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n393), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  AND2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(G1333gat));
  XNOR2_X1  g559(.A(new_n516), .B(KEYINPUT107), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n750), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n695), .A2(G71gat), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n762), .A2(G71gat), .B1(new_n752), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g564(.A1(new_n679), .A2(new_n422), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT108), .B(G78gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n562), .A2(new_n648), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n748), .A2(new_n703), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n770), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n714), .B2(new_n523), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n703), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n679), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n286), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n574), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n770), .A2(new_n751), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n710), .B2(new_n722), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(new_n286), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(KEYINPUT109), .A3(new_n778), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n779), .B1(new_n786), .B2(new_n574), .ZN(G1336gat));
  NOR3_X1   g586(.A1(new_n679), .A2(G92gat), .A3(new_n393), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n771), .A2(new_n772), .ZN(new_n789));
  XNOR2_X1  g588(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n775), .B2(new_n703), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(KEYINPUT111), .B(new_n788), .C1(new_n789), .C2(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n289), .B1(new_n782), .B2(new_n504), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n797), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n393), .A2(G92gat), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(new_n777), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(G1337gat));
  XNOR2_X1  g602(.A(KEYINPUT112), .B(G99gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n777), .A2(new_n697), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n695), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n783), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n807), .B2(new_n804), .ZN(G1338gat));
  AOI21_X1  g607(.A(new_n414), .B1(new_n782), .B2(new_n423), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n789), .A2(new_n791), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n766), .A2(new_n414), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT113), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n782), .B2(new_n423), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n709), .A2(KEYINPUT44), .B1(new_n721), .B2(new_n715), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n817), .A2(KEYINPUT114), .A3(new_n422), .A4(new_n781), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n816), .A2(new_n818), .A3(new_n414), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n773), .A2(new_n776), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n811), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n814), .B1(new_n819), .B2(new_n822), .ZN(G1339gat));
  NOR3_X1   g622(.A1(new_n622), .A2(new_n648), .A3(new_n751), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n658), .A2(new_n665), .A3(new_n659), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n827));
  AOI21_X1  g626(.A(new_n671), .B1(new_n673), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT55), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  INV_X1    g629(.A(new_n672), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n626), .B1(new_n625), .B2(new_n628), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n634), .B1(new_n633), .B2(new_n636), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n643), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n647), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n832), .A2(new_n719), .A3(new_n720), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n832), .A2(new_n648), .B1(new_n751), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n721), .ZN(new_n840));
  INV_X1    g639(.A(new_n562), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n824), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n753), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n510), .A2(new_n513), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT117), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n393), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT118), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n849), .A3(new_n393), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n648), .A2(new_n205), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT119), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n842), .B2(new_n423), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n646), .A2(new_n647), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n826), .A2(new_n828), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n672), .A3(new_n860), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n856), .A2(new_n861), .B1(new_n679), .B2(new_n836), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n719), .A2(new_n720), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n562), .B1(new_n864), .B2(new_n838), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n855), .B(new_n422), .C1(new_n865), .C2(new_n824), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n854), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n286), .A2(new_n504), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n697), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n856), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n870), .ZN(G1340gat));
  NAND2_X1  g670(.A1(new_n751), .A2(new_n203), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT120), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n848), .A2(new_n850), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G120gat), .B1(new_n869), .B2(new_n679), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1341gat));
  NOR3_X1   g675(.A1(new_n869), .A2(new_n211), .A3(new_n841), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n846), .A2(new_n393), .A3(new_n562), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n211), .ZN(G1342gat));
  NOR2_X1   g678(.A1(new_n621), .A2(G134gat), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n847), .A2(KEYINPUT56), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n869), .B2(new_n621), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT56), .B1(new_n847), .B2(new_n881), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1343gat));
  INV_X1    g684(.A(new_n842), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n423), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n806), .A2(new_n868), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n857), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT55), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n830), .A2(new_n891), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n648), .A3(new_n672), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n751), .A2(new_n837), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n703), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n838), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n841), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n824), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n422), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n888), .B(new_n890), .C1(new_n887), .C2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G141gat), .B1(new_n902), .B2(new_n856), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n695), .A2(new_n422), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n843), .A2(new_n393), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n218), .A3(new_n648), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n220), .A3(new_n751), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n887), .B1(new_n886), .B2(new_n423), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n861), .A2(new_n621), .A3(new_n836), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n841), .B1(new_n897), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n900), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n422), .A2(KEYINPUT57), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n889), .A2(KEYINPUT122), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n889), .A2(KEYINPUT122), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n916), .A2(new_n751), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n910), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n910), .B(G148gat), .C1(new_n902), .C2(new_n679), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n909), .B1(new_n920), .B2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(G155gat), .B1(new_n905), .B2(new_n562), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n902), .A2(new_n224), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n562), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n902), .B2(new_n863), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n225), .A3(new_n703), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n842), .A2(new_n778), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n844), .A2(new_n504), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT123), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n310), .A3(new_n648), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n753), .A2(new_n504), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n867), .A2(new_n761), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(new_n648), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n937), .B2(new_n310), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n936), .A2(G176gat), .A3(new_n751), .ZN(new_n939));
  INV_X1    g738(.A(new_n933), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n311), .B1(new_n940), .B2(new_n679), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(G1349gat));
  AOI21_X1  g741(.A(new_n337), .B1(new_n936), .B2(new_n562), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n933), .A2(new_n359), .A3(new_n562), .ZN(new_n944));
  OR3_X1    g743(.A1(new_n943), .A2(KEYINPUT60), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT60), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n933), .A2(new_n358), .A3(new_n721), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n867), .A2(new_n703), .A3(new_n761), .A4(new_n935), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n949), .A2(new_n950), .A3(G190gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n949), .B2(G190gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(new_n948), .C1(new_n951), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1351gat));
  NAND3_X1  g756(.A1(new_n930), .A2(new_n504), .A3(new_n904), .ZN(new_n958));
  XNOR2_X1  g757(.A(KEYINPUT125), .B(G197gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n958), .A2(new_n856), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n935), .A2(new_n806), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n916), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n959), .B1(new_n964), .B2(new_n856), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n961), .A2(new_n965), .ZN(G1352gat));
  INV_X1    g765(.A(new_n958), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(new_n669), .A3(new_n751), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n916), .A2(new_n751), .A3(new_n963), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G204gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n968), .B2(KEYINPUT62), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n970), .A2(new_n971), .A3(new_n973), .A4(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n967), .A2(new_n292), .A3(new_n562), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n916), .A2(new_n562), .A3(new_n963), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n964), .B2(new_n621), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n967), .A2(new_n293), .A3(new_n721), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


