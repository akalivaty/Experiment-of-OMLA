//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(KEYINPUT84), .B(G29gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(G36gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT14), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G43gat), .B(G50gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT83), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT83), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(KEYINPUT15), .A3(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT85), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n202), .A2(G36gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n205), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(KEYINPUT85), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n216), .A2(new_n212), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n213), .A2(KEYINPUT17), .A3(new_n219), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G1gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n225), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G8gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(new_n229), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n233), .A3(new_n230), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n220), .B(new_n229), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n236), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT82), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT11), .B(G169gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n242), .B(new_n245), .C1(KEYINPUT87), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT87), .A3(new_n241), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n243), .A2(new_n244), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n241), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(G85gat), .A2(G92gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT7), .ZN(new_n261));
  XNOR2_X1  g060(.A(G99gat), .B(G106gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263));
  INV_X1    g062(.A(G85gat), .ZN(new_n264));
  INV_X1    g063(.A(G92gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(KEYINPUT8), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n262), .B1(new_n261), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT98), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT98), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT89), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(G71gat), .A2(G78gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT9), .ZN(new_n278));
  INV_X1    g077(.A(G71gat), .ZN(new_n279));
  INV_X1    g078(.A(G78gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n277), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT9), .ZN(new_n285));
  OAI221_X1 g084(.A(new_n284), .B1(new_n285), .B2(new_n274), .C1(new_n279), .C2(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT90), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n286), .A3(KEYINPUT90), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n289), .A2(KEYINPUT95), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT95), .B1(new_n289), .B2(new_n290), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT10), .B(new_n273), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT10), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n269), .A2(new_n282), .A3(new_n286), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n290), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n294), .B(new_n295), .C1(new_n297), .C2(new_n273), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n259), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n273), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n259), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(G204gat), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n301), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n258), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT65), .B(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT27), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n313));
  INV_X1    g112(.A(G190gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT27), .B(G183gat), .Z(new_n316));
  OAI21_X1  g115(.A(KEYINPUT28), .B1(new_n316), .B2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  OR3_X1    g117(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(G169gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(new_n303), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n315), .A2(new_n317), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n321), .A3(new_n303), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  AOI211_X1 g129(.A(new_n330), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G183gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n314), .ZN(new_n336));
  NAND3_X1  g135(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT25), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(KEYINPUT65), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  AOI21_X1  g141(.A(G190gat), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n337), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n328), .B(KEYINPUT25), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT66), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n334), .B(new_n337), .C1(new_n309), .C2(G190gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT25), .A4(new_n328), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n323), .B1(new_n339), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(G120gat), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n358));
  INV_X1    g157(.A(G120gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G134gat), .ZN(new_n363));
  INV_X1    g162(.A(G134gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G127gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n365), .A3(KEYINPUT67), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367));
  NAND2_X1  g166(.A1(G113gat), .A2(G120gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n360), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OR3_X1    g168(.A1(new_n364), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n361), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n351), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n338), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n329), .A2(new_n331), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n346), .B(new_n349), .C1(new_n375), .C2(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n371), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n323), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n373), .A2(G227gat), .A3(G233gat), .A4(new_n378), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT34), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT32), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n383), .B2(KEYINPUT32), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(KEYINPUT32), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n385), .A3(new_n381), .ZN(new_n391));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G71gat), .ZN(new_n393));
  INV_X1    g192(.A(G99gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n383), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(KEYINPUT33), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n388), .A2(new_n391), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n388), .B2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT36), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n386), .A2(new_n387), .A3(new_n382), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n381), .B1(new_n390), .B2(new_n385), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n397), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT36), .B1(new_n406), .B2(new_n399), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT28), .B(G190gat), .C1(new_n310), .C2(new_n311), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n317), .A2(new_n318), .A3(new_n322), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n346), .A2(new_n349), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n338), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n412), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n409), .B1(new_n419), .B2(KEYINPUT29), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT71), .B1(new_n419), .B2(new_n409), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT71), .ZN(new_n422));
  INV_X1    g221(.A(new_n409), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n351), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT22), .ZN(new_n427));
  INV_X1    g226(.A(G211gat), .ZN(new_n428));
  INV_X1    g227(.A(G218gat), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G211gat), .B(G218gat), .Z(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT70), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n434), .A2(new_n435), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n425), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT37), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n351), .A2(new_n423), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT29), .B1(new_n376), .B2(new_n323), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n441), .B(new_n437), .C1(new_n442), .C2(new_n423), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT72), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT72), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n420), .A2(new_n445), .A3(new_n437), .A4(new_n441), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n439), .A2(new_n440), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448));
  INV_X1    g247(.A(G64gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(new_n265), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n439), .A2(new_n444), .A3(new_n446), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(KEYINPUT37), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n447), .B1(new_n454), .B2(KEYINPUT81), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  AOI211_X1 g255(.A(new_n456), .B(new_n452), .C1(new_n453), .C2(KEYINPUT37), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT38), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G141gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(G148gat), .ZN(new_n460));
  INV_X1    g259(.A(G148gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(G141gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT74), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(G141gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(G148gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT74), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n463), .A2(new_n464), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G155gat), .B(G162gat), .Z(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OR3_X1    g271(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n473), .A2(new_n474), .B1(new_n465), .B2(new_n466), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n372), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT4), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT77), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n470), .B2(new_n471), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n372), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n472), .A2(new_n476), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT3), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n377), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n361), .A2(new_n371), .A3(KEYINPUT76), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n480), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n486), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n483), .A2(new_n484), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT78), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g297(.A(new_n490), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n477), .B1(new_n499), .B2(new_n480), .ZN(new_n500));
  INV_X1    g299(.A(new_n484), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n491), .B1(new_n472), .B2(new_n476), .ZN(new_n503));
  AOI211_X1 g302(.A(KEYINPUT3), .B(new_n475), .C1(new_n470), .C2(new_n471), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n505), .B2(new_n490), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(KEYINPUT78), .A3(new_n483), .A4(new_n494), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n497), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G1gat), .B(G29gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT0), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G57gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(new_n264), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n478), .A2(new_n482), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n498), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n508), .B2(new_n514), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n508), .A2(new_n514), .ZN(new_n520));
  INV_X1    g319(.A(new_n512), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT6), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n425), .A2(new_n437), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n420), .A2(new_n438), .A3(new_n441), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT37), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT38), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n447), .A2(new_n527), .A3(new_n528), .A4(new_n451), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n439), .A2(new_n444), .A3(new_n446), .A4(new_n452), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n458), .A2(new_n524), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G50gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G228gat), .A2(G233gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n434), .A2(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n432), .A2(new_n433), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT3), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n538), .B2(new_n480), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n437), .B1(new_n492), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n437), .A2(new_n540), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n480), .B1(new_n543), .B2(new_n491), .ZN(new_n544));
  OAI211_X1 g343(.A(G228gat), .B(G233gat), .C1(new_n544), .C2(new_n541), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n534), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G78gat), .B(G106gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G22gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT79), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n542), .A2(new_n545), .A3(new_n534), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n550), .ZN(new_n553));
  INV_X1    g352(.A(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n444), .A2(new_n446), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT71), .B(new_n409), .C1(new_n376), .C2(new_n323), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n422), .B1(new_n351), .B2(new_n423), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n437), .B1(new_n560), .B2(new_n420), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n562), .A2(KEYINPUT73), .A3(KEYINPUT30), .A4(new_n452), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n530), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n451), .B1(new_n557), .B2(new_n561), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT30), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n530), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT39), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n484), .B1(new_n513), .B2(new_n493), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT80), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(KEYINPUT80), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n573), .A2(KEYINPUT80), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n500), .A2(new_n501), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(new_n572), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n512), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n520), .A2(new_n521), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n577), .A2(new_n581), .A3(KEYINPUT40), .A4(new_n512), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n556), .B1(new_n571), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n408), .B1(new_n532), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n516), .A3(new_n515), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n522), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(new_n570), .A3(new_n567), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n556), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595));
  INV_X1    g394(.A(new_n556), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n406), .A3(new_n399), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n400), .A2(new_n556), .A3(new_n401), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n566), .A2(new_n563), .B1(new_n569), .B2(new_n530), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(KEYINPUT35), .A3(new_n591), .A4(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  INV_X1    g405(.A(new_n292), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n289), .A2(KEYINPUT95), .A3(new_n290), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n605), .B1(new_n609), .B2(new_n229), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT21), .B1(new_n291), .B2(new_n292), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n230), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n610), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n604), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT94), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n616), .B2(new_n620), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n296), .A2(new_n606), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT19), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n622), .B2(new_n623), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n270), .A2(KEYINPUT99), .A3(new_n272), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n222), .A3(new_n223), .ZN(new_n639));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n213), .B(new_n219), .C1(KEYINPUT99), .C2(KEYINPUT17), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n273), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n314), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n314), .B1(new_n639), .B2(new_n644), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n429), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(G218gat), .A3(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n640), .A2(new_n641), .ZN(new_n655));
  INV_X1    g454(.A(G162gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT97), .B(G134gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n652), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n654), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n308), .A2(new_n603), .A3(new_n637), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n524), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n571), .ZN(new_n666));
  NOR2_X1   g465(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n667));
  AND2_X1   g466(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n666), .A2(G8gat), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT42), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(KEYINPUT42), .B2(new_n669), .ZN(G1325gat));
  NOR2_X1   g471(.A1(new_n400), .A2(new_n401), .ZN(new_n673));
  AOI21_X1  g472(.A(G15gat), .B1(new_n663), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n408), .A2(G15gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n663), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n663), .A2(new_n556), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  AOI21_X1  g478(.A(new_n662), .B1(new_n594), .B2(new_n602), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n634), .A2(new_n636), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(new_n308), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n683), .A2(new_n591), .A3(new_n202), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT45), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n598), .A2(new_n601), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n689), .B(new_n596), .C1(new_n600), .C2(new_n591), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT101), .B1(new_n592), .B2(new_n556), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n688), .B1(new_n692), .B2(new_n589), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n687), .B1(new_n693), .B2(new_n662), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n686), .A2(new_n694), .A3(new_n682), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n202), .B1(new_n695), .B2(new_n591), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n685), .A2(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n683), .A2(G36gat), .A3(new_n600), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n695), .B2(new_n600), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n673), .A2(KEYINPUT36), .ZN(new_n702));
  INV_X1    g501(.A(new_n407), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G43gat), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n673), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n683), .A2(G43gat), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT47), .B1(new_n707), .B2(KEYINPUT102), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1330gat));
  INV_X1    g509(.A(G50gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n683), .B2(new_n596), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n596), .A2(new_n711), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n686), .A2(new_n694), .A3(new_n682), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT103), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g516(.A(new_n258), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n693), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n662), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n681), .A2(new_n306), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n591), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT104), .B(G57gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1332gat));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n571), .B1(new_n726), .B2(new_n449), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT105), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n719), .A2(new_n721), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n449), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1333gat));
  OAI21_X1  g530(.A(new_n279), .B1(new_n722), .B2(new_n706), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n408), .A2(G71gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n722), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n722), .A2(new_n596), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n280), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n637), .A2(new_n718), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n686), .A2(new_n694), .A3(new_n307), .A4(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n264), .A3(new_n591), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n693), .B2(new_n662), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n593), .A2(new_n689), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n592), .A2(KEYINPUT101), .A3(new_n556), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n590), .A2(new_n522), .A3(new_n530), .A4(new_n529), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n451), .B1(new_n562), .B2(new_n440), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n456), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n447), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(KEYINPUT38), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n596), .B1(new_n600), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n704), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n602), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n720), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n756), .A3(new_n738), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n756), .A3(KEYINPUT51), .A4(new_n738), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n306), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n524), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n740), .B1(new_n762), .B2(new_n264), .ZN(G1336gat));
  NOR3_X1   g562(.A1(new_n739), .A2(new_n265), .A3(new_n600), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n759), .A2(new_n760), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n307), .A3(new_n571), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(new_n766), .B2(new_n265), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT52), .B1(new_n767), .B2(KEYINPUT107), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  AOI21_X1  g569(.A(G92gat), .B1(new_n761), .B2(new_n571), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n764), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1337gat));
  AOI21_X1  g572(.A(G99gat), .B1(new_n761), .B2(new_n673), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n739), .A2(new_n394), .A3(new_n704), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1338gat));
  XOR2_X1   g578(.A(KEYINPUT109), .B(G106gat), .Z(new_n780));
  OAI211_X1 g579(.A(KEYINPUT110), .B(new_n780), .C1(new_n739), .C2(new_n596), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n306), .A2(G106gat), .A3(new_n596), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT111), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n759), .B2(new_n760), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT53), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n780), .B1(new_n739), .B2(new_n596), .ZN(new_n788));
  NAND2_X1  g587(.A1(KEYINPUT110), .A2(KEYINPUT53), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n759), .B2(new_n760), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n787), .B(KEYINPUT112), .C1(new_n790), .C2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n784), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n791), .B1(new_n796), .B2(new_n781), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n790), .A2(new_n793), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(G1339gat));
  AND3_X1   g599(.A1(new_n306), .A2(new_n253), .A3(new_n257), .ZN(new_n801));
  AND4_X1   g600(.A1(new_n634), .A2(new_n636), .A3(new_n662), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n236), .B1(new_n235), .B2(new_n237), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n239), .A2(new_n240), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n250), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n242), .A2(new_n252), .A3(new_n245), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n662), .A2(new_n307), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n258), .A2(new_n662), .ZN(new_n808));
  INV_X1    g607(.A(new_n305), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n301), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n299), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n305), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n815), .A3(new_n305), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n293), .A2(new_n259), .A3(new_n298), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n819), .A2(new_n299), .A3(new_n811), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT55), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n815), .B1(new_n812), .B2(new_n305), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT113), .B(new_n809), .C1(new_n299), .C2(new_n811), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT55), .B(new_n820), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n806), .A2(new_n805), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n660), .A3(new_n661), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n808), .A2(new_n810), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n817), .A2(new_n820), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT55), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n807), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n802), .B1(new_n832), .B2(new_n681), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n591), .A3(new_n571), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n599), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n258), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n354), .A2(new_n355), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n353), .B2(new_n836), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n835), .A2(new_n306), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(new_n359), .ZN(G1341gat));
  NOR2_X1   g640(.A1(new_n835), .A2(new_n681), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G127gat), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n842), .A2(G127gat), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1342gat));
  AOI211_X1 g646(.A(new_n662), .B(new_n835), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT116), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n848), .B(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT58), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n833), .B2(new_n596), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n828), .A2(new_n810), .ZN(new_n857));
  INV_X1    g656(.A(new_n831), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n808), .A4(new_n826), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n637), .B1(new_n859), .B2(new_n807), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT57), .B(new_n556), .C1(new_n860), .C2(new_n802), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT117), .B(new_n854), .C1(new_n833), .C2(new_n596), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n571), .A2(new_n591), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n704), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n718), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n852), .A2(KEYINPUT58), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n408), .A2(new_n596), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n834), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n718), .A2(new_n459), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT118), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n853), .A2(new_n868), .A3(new_n869), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n867), .B2(G141gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n853), .B1(new_n877), .B2(new_n869), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(new_n871), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n461), .A3(new_n307), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n307), .A2(new_n862), .A3(new_n863), .A4(new_n866), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(KEYINPUT59), .A3(new_n461), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n855), .A2(new_n861), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n307), .A3(new_n866), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n881), .B1(new_n883), .B2(new_n887), .ZN(G1345gat));
  INV_X1    g687(.A(G155gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n889), .A3(new_n637), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n637), .A2(new_n862), .A3(new_n863), .A4(new_n866), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n889), .ZN(G1346gat));
  NAND3_X1  g691(.A1(new_n880), .A2(new_n656), .A3(new_n720), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n720), .A2(new_n862), .A3(new_n863), .A4(new_n866), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n656), .ZN(G1347gat));
  OAI21_X1  g694(.A(KEYINPUT121), .B1(new_n833), .B2(new_n524), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n597), .A2(new_n600), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n898), .B(new_n591), .C1(new_n860), .C2(new_n802), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT122), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n321), .A3(new_n718), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n897), .B(new_n591), .C1(new_n860), .C2(new_n802), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n258), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1348gat));
  NOR3_X1   g704(.A1(new_n903), .A2(new_n303), .A3(new_n306), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n901), .A2(new_n307), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n303), .ZN(G1349gat));
  NOR2_X1   g707(.A1(new_n681), .A2(new_n316), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n896), .A2(new_n899), .A3(new_n897), .A4(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n309), .B1(new_n903), .B2(new_n681), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT123), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n314), .A3(new_n720), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n903), .B2(new_n662), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n408), .A2(new_n600), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n591), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT125), .Z(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n885), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n258), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n896), .A2(new_n899), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n556), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT124), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n258), .A2(G197gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  XNOR2_X1  g733(.A(KEYINPUT126), .B(G204gat), .ZN(new_n935));
  OR4_X1    g734(.A1(KEYINPUT62), .A2(new_n932), .A3(new_n306), .A4(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n885), .A2(new_n307), .A3(new_n925), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n935), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n929), .A2(new_n931), .ZN(new_n939));
  INV_X1    g738(.A(new_n935), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n307), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n938), .A3(new_n942), .ZN(G1353gat));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n681), .B(new_n924), .C1(new_n855), .C2(new_n861), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n428), .ZN(new_n946));
  OAI211_X1 g745(.A(KEYINPUT63), .B(G211gat), .C1(new_n926), .C2(new_n681), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT127), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n939), .A2(new_n428), .A3(new_n637), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n950), .B(new_n944), .C1(new_n945), .C2(new_n428), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(G1354gat));
  NOR3_X1   g751(.A1(new_n926), .A2(new_n429), .A3(new_n662), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n939), .A2(new_n720), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n429), .ZN(G1355gat));
endmodule


