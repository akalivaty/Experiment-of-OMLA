//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202));
  INV_X1    g001(.A(G230gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  OR2_X1    g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT96), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G64gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n213), .A2(G57gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(G57gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT9), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n216), .A2(KEYINPUT96), .A3(new_n206), .A4(new_n207), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n206), .B1(new_n207), .B2(new_n209), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n214), .B2(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT7), .ZN(new_n222));
  INV_X1    g021(.A(G99gat), .ZN(new_n223));
  INV_X1    g022(.A(G106gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT8), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G85gat), .ZN(new_n226));
  INV_X1    g025(.A(G92gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n225), .A2(KEYINPUT98), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT98), .B1(new_n225), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n222), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G99gat), .B(G106gat), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n232), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n222), .C1(new_n229), .C2(new_n230), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n220), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT10), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n235), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n212), .A2(new_n220), .A3(new_n217), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n236), .A3(new_n237), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n205), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n205), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(new_n241), .B2(new_n236), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n202), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G120gat), .B(G148gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(G176gat), .B(G204gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n246), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT23), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n254), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n255), .B2(new_n252), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT25), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G183gat), .ZN(new_n262));
  INV_X1    g061(.A(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n259), .A2(KEYINPUT64), .A3(KEYINPUT24), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT24), .B1(new_n259), .B2(KEYINPUT64), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n269), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n256), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n261), .B1(new_n271), .B2(KEYINPUT25), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G183gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT27), .B(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n273), .B1(new_n282), .B2(new_n263), .ZN(new_n283));
  INV_X1    g082(.A(new_n259), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n274), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n286), .B(new_n263), .C1(new_n285), .C2(new_n279), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n252), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n283), .A2(new_n284), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n296));
  OAI21_X1  g095(.A(G134gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(KEYINPUT70), .B(G134gat), .C1(new_n295), .C2(new_n296), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n301), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT68), .B1(new_n301), .B2(G127gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G120gat), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G113gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT71), .B1(new_n309), .B2(G113gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(new_n307), .A3(G120gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n316), .C1(new_n307), .C2(G120gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n306), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n312), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n313), .B1(new_n312), .B2(new_n319), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n272), .A2(new_n294), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n259), .A2(KEYINPUT64), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n259), .A2(KEYINPUT64), .A3(KEYINPUT24), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n269), .B1(new_n327), .B2(new_n264), .ZN(new_n328));
  INV_X1    g127(.A(new_n270), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT25), .B(new_n257), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n261), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n319), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n312), .A2(new_n313), .A3(new_n319), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n278), .A2(new_n281), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT28), .B1(new_n336), .B2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n293), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n259), .A3(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT34), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n342), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n340), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350));
  INV_X1    g149(.A(G43gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT73), .B(G15gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT33), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n349), .A2(KEYINPUT32), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n349), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n349), .A2(KEYINPUT32), .ZN(new_n361));
  INV_X1    g160(.A(new_n349), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n361), .B(new_n354), .C1(new_n362), .C2(KEYINPUT33), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n347), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n363), .ZN(new_n365));
  INV_X1    g164(.A(new_n346), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n345), .B(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n370), .B(KEYINPUT86), .Z(new_n371));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n372));
  INV_X1    g171(.A(G141gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(G148gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(G148gat), .ZN(new_n375));
  INV_X1    g174(.A(G148gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT79), .A3(G141gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G155gat), .B(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT2), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G155gat), .B(G162gat), .Z(new_n383));
  XNOR2_X1  g182(.A(G141gat), .B(G148gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(KEYINPUT2), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387));
  INV_X1    g186(.A(G211gat), .ZN(new_n388));
  INV_X1    g187(.A(G218gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT22), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT87), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(KEYINPUT22), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n387), .A3(new_n390), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n386), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n394), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n385), .A3(new_n401), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n371), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n382), .A2(new_n385), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(KEYINPUT88), .A3(new_n399), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n401), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT88), .B1(new_n403), .B2(new_n399), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n405), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n411), .A2(G228gat), .A3(G233gat), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT31), .B(G50gat), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G22gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n416), .B(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n369), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT35), .ZN(new_n422));
  INV_X1    g221(.A(new_n403), .ZN(new_n423));
  INV_X1    g222(.A(G226gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(new_n204), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n272), .A2(new_n294), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(KEYINPUT29), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n332), .B2(new_n339), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(new_n227), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT77), .B(G64gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI22_X1  g233(.A1(new_n272), .A2(new_n294), .B1(KEYINPUT29), .B2(new_n425), .ZN(new_n435));
  INV_X1    g234(.A(new_n425), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n332), .A2(new_n339), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n437), .A3(new_n403), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n439), .A2(KEYINPUT78), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n439), .B2(KEYINPUT78), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n429), .B2(new_n438), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT82), .B(G1gat), .Z(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n447), .B(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n317), .A2(new_n306), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n452), .A2(new_n318), .B1(new_n305), .B2(new_n311), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n386), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n333), .A2(new_n407), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT4), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n407), .A2(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n404), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n463), .B2(new_n453), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n464), .A2(new_n454), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT4), .B(new_n386), .C1(new_n320), .C2(new_n321), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n459), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n312), .A2(new_n386), .A3(new_n319), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n382), .A2(new_n385), .A3(new_n401), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n401), .B1(new_n382), .B2(new_n385), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n469), .A2(KEYINPUT4), .B1(new_n472), .B2(new_n333), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n407), .B1(new_n334), .B2(new_n335), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(KEYINPUT4), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n450), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n475), .A2(KEYINPUT4), .B1(new_n454), .B2(new_n464), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n386), .B1(new_n312), .B2(new_n319), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n469), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT5), .B1(new_n482), .B2(new_n457), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n476), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n486), .A3(new_n476), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n450), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n478), .ZN(new_n489));
  INV_X1    g288(.A(new_n450), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n479), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n421), .A2(new_n422), .A3(new_n444), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n416), .B(new_n418), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n368), .B2(new_n364), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT84), .B1(new_n491), .B2(new_n477), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n484), .A2(new_n490), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n468), .A2(new_n476), .A3(new_n450), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n489), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n479), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n501), .A2(new_n502), .A3(new_n444), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n501), .B2(new_n444), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n495), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n493), .B1(new_n505), .B2(new_n422), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n312), .A2(new_n386), .A3(KEYINPUT4), .A4(new_n319), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n463), .B2(new_n453), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n386), .B1(new_n320), .B2(new_n321), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(new_n460), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n511), .A2(new_n512), .A3(new_n457), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n473), .B1(new_n475), .B2(KEYINPUT4), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT89), .B1(new_n514), .B2(new_n458), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n507), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n512), .B1(new_n511), .B2(new_n457), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n334), .A2(new_n335), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT4), .B1(new_n518), .B2(new_n386), .ZN(new_n519));
  OAI211_X1 g318(.A(KEYINPUT89), .B(new_n458), .C1(new_n519), .C2(new_n509), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n507), .B1(new_n482), .B2(new_n457), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n450), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT90), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n488), .B1(new_n524), .B2(KEYINPUT40), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n517), .A2(new_n520), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n490), .B1(new_n527), .B2(new_n507), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n444), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n420), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533));
  INV_X1    g332(.A(new_n438), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n403), .B1(new_n435), .B2(new_n437), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT37), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT38), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT37), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n429), .A2(new_n538), .A3(new_n438), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n433), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n439), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n533), .B1(new_n492), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n433), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT38), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n486), .B1(new_n468), .B2(new_n476), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n490), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n491), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n540), .A2(new_n439), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT92), .A4(new_n479), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n542), .A2(new_n544), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n420), .B1(new_n503), .B2(new_n504), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n365), .A2(new_n367), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n347), .A2(new_n360), .A3(new_n363), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT76), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT36), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n251), .B1(new_n506), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G197gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT11), .B(G169gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT12), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n567));
  INV_X1    g366(.A(G29gat), .ZN(new_n568));
  INV_X1    g367(.A(G36gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n570), .A2(new_n571), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n351), .A2(G50gat), .ZN(new_n574));
  INV_X1    g373(.A(G50gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(G43gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n573), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G43gat), .B(G50gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT15), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n572), .A2(new_n581), .A3(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(G15gat), .A2(G22gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g384(.A1(G15gat), .A2(G22gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n588), .A2(G1gat), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT16), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(G1gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT94), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n594), .B2(new_n587), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n590), .A2(new_n595), .A3(G8gat), .ZN(new_n596));
  INV_X1    g395(.A(G8gat), .ZN(new_n597));
  OAI22_X1  g396(.A1(new_n588), .A2(new_n589), .B1(new_n591), .B2(G1gat), .ZN(new_n598));
  INV_X1    g397(.A(G1gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n599), .A3(new_n587), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n583), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(G8gat), .B1(new_n590), .B2(new_n595), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n597), .A3(new_n600), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n580), .A4(new_n582), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT13), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT95), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n580), .A2(KEYINPUT17), .A3(new_n582), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(new_n582), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n581), .B1(new_n577), .B2(new_n572), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n613), .A2(new_n617), .A3(new_n603), .A4(new_n604), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n602), .ZN(new_n619));
  INV_X1    g418(.A(new_n607), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT18), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n618), .A2(new_n602), .A3(new_n622), .A4(new_n607), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n610), .A2(new_n612), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n566), .B1(new_n625), .B2(KEYINPUT93), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n624), .A2(new_n627), .A3(new_n565), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n560), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT97), .Z(new_n633));
  NAND4_X1  g432(.A1(new_n212), .A2(new_n217), .A3(KEYINPUT21), .A4(new_n220), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n603), .A2(new_n634), .A3(new_n604), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G183gat), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n603), .A2(new_n634), .A3(new_n604), .A4(new_n262), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n633), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n637), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n638), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n645));
  INV_X1    g444(.A(new_n633), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n240), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n388), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n649), .B(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n642), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n642), .B2(new_n647), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G134gat), .B(G162gat), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n239), .A2(new_n613), .A3(new_n617), .ZN(new_n659));
  XOR2_X1   g458(.A(G190gat), .B(G218gat), .Z(new_n660));
  NAND3_X1  g459(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n583), .A2(new_n235), .A3(new_n233), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n658), .B1(new_n664), .B2(KEYINPUT99), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n666));
  INV_X1    g465(.A(new_n660), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n669), .A3(new_n663), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n658), .A3(new_n663), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n668), .A2(KEYINPUT100), .A3(new_n658), .A4(new_n663), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n642), .A2(new_n647), .ZN(new_n679));
  INV_X1    g478(.A(new_n652), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n642), .A2(new_n647), .A3(new_n652), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n678), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n631), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n501), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT103), .B(G1gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1324gat));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n444), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(KEYINPUT42), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(KEYINPUT105), .B2(new_n693), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(KEYINPUT105), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n691), .A2(new_n597), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n694), .B1(new_n696), .B2(new_n699), .ZN(G1325gat));
  NOR2_X1   g499(.A1(new_n687), .A2(new_n369), .ZN(new_n701));
  INV_X1    g500(.A(new_n558), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G15gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT106), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI22_X1  g504(.A1(new_n701), .A2(G15gat), .B1(new_n687), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT107), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n687), .A2(new_n494), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NAND3_X1  g509(.A1(new_n560), .A2(new_n655), .A3(new_n630), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n684), .ZN(new_n712));
  INV_X1    g511(.A(new_n501), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n568), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n559), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n553), .A2(new_n558), .A3(new_n554), .A4(KEYINPUT109), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n506), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n719), .B2(new_n676), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n506), .A2(new_n559), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n721), .A2(KEYINPUT44), .A3(new_n676), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n250), .B(KEYINPUT108), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n683), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n720), .A2(new_n722), .A3(new_n629), .A4(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n713), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n715), .B1(new_n568), .B2(new_n728), .ZN(G1328gat));
  INV_X1    g528(.A(new_n712), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(G36gat), .A3(new_n444), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g533(.A(new_n444), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n733), .B(new_n734), .C1(new_n569), .C2(new_n736), .ZN(G1329gat));
  NOR4_X1   g536(.A1(new_n711), .A2(G43gat), .A3(new_n684), .A4(new_n369), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n720), .A2(new_n722), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n739), .A2(new_n630), .A3(new_n702), .A4(new_n725), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT47), .B(new_n738), .C1(new_n740), .C2(G43gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(G1330gat));
  NOR3_X1   g544(.A1(new_n730), .A2(G50gat), .A3(new_n494), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n727), .A2(new_n420), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n575), .ZN(new_n750));
  INV_X1    g549(.A(new_n748), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n575), .B1(new_n727), .B2(new_n420), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n746), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(G1331gat));
  NOR3_X1   g553(.A1(new_n630), .A2(new_n677), .A3(new_n685), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n719), .A2(new_n724), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n719), .A2(new_n758), .A3(new_n724), .A4(new_n755), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n713), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n735), .A3(new_n759), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT49), .B(G64gat), .Z(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(G1333gat));
  NAND3_X1  g564(.A1(new_n757), .A2(new_n702), .A3(new_n759), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G71gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n369), .A2(G71gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n757), .A2(new_n759), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1334gat));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n420), .A3(new_n759), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n630), .A2(new_n683), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n251), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n720), .A2(new_n722), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n501), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n719), .A2(new_n676), .A3(new_n775), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n719), .A2(KEYINPUT51), .A3(new_n676), .A4(new_n775), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(new_n226), .A3(new_n713), .A4(new_n251), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n785), .ZN(G1336gat));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n227), .B1(new_n777), .B2(new_n735), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n735), .A2(new_n227), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n723), .B(new_n789), .C1(new_n782), .C2(new_n783), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT112), .B(new_n787), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n784), .A2(new_n227), .A3(new_n735), .A4(new_n724), .ZN(new_n792));
  INV_X1    g591(.A(new_n720), .ZN(new_n793));
  INV_X1    g592(.A(new_n722), .ZN(new_n794));
  INV_X1    g593(.A(new_n776), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n793), .A2(new_n735), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n791), .A2(new_n800), .ZN(G1337gat));
  XOR2_X1   g600(.A(KEYINPUT113), .B(G99gat), .Z(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n778), .B2(new_n558), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n369), .A2(new_n802), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n251), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1338gat));
  NOR2_X1   g605(.A1(new_n494), .A2(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n784), .A2(new_n724), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n224), .B1(new_n777), .B2(new_n420), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n810), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n808), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n686), .A2(new_n816), .A3(new_n629), .A4(new_n250), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT101), .B1(new_n655), .B2(new_n676), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n683), .A2(new_n684), .A3(new_n678), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n629), .A3(new_n819), .A4(new_n250), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n606), .A2(new_n608), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n619), .A2(new_n620), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n564), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n624), .B2(new_n565), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n676), .B1(new_n251), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT115), .A4(new_n205), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n238), .A2(new_n242), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n244), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n244), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT54), .B(new_n827), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n249), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n243), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n243), .A2(new_n245), .A3(new_n249), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n826), .B1(new_n841), .B2(new_n629), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n838), .A2(new_n825), .A3(new_n839), .A4(new_n840), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n683), .B1(new_n843), .B2(new_n676), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n817), .A2(new_n821), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n495), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n501), .A2(new_n735), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n629), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT116), .B(G113gat), .Z(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n848), .B2(new_n723), .ZN(new_n852));
  INV_X1    g651(.A(new_n847), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n250), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n846), .A2(new_n309), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(G1341gat));
  INV_X1    g655(.A(new_n848), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n683), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n295), .A2(new_n296), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(G1342gat));
  NOR2_X1   g659(.A1(new_n848), .A2(new_n684), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n301), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT117), .ZN(new_n864));
  INV_X1    g663(.A(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G134gat), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT56), .B1(new_n865), .B2(G134gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n864), .A2(KEYINPUT118), .A3(new_n866), .A4(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1343gat));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n845), .A2(new_n873), .A3(new_n494), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n853), .B1(new_n874), .B2(KEYINPUT119), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n817), .A2(new_n821), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n844), .A2(new_n842), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .A3(new_n420), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n845), .B2(new_n494), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n558), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G141gat), .B1(new_n883), .B2(new_n629), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n845), .A2(new_n702), .A3(new_n494), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n847), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n630), .A2(new_n373), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n702), .B1(new_n874), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n877), .A2(new_n820), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n873), .B1(new_n894), .B2(new_n494), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n879), .A3(KEYINPUT121), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n896), .A3(new_n854), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n891), .B1(new_n897), .B2(G148gat), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n875), .A2(new_n882), .A3(new_n558), .A4(new_n251), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n376), .A2(KEYINPUT59), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT120), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n899), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n898), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n886), .A2(G148gat), .A3(new_n250), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n890), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n906), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n899), .A2(new_n903), .A3(new_n900), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n899), .B2(new_n900), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT122), .B(new_n908), .C1(new_n911), .C2(new_n898), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n907), .A2(new_n912), .ZN(G1345gat));
  XNOR2_X1  g712(.A(KEYINPUT80), .B(G155gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n883), .A2(new_n655), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n885), .A2(new_n683), .A3(new_n847), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(G1346gat));
  INV_X1    g717(.A(G162gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n883), .A2(new_n919), .A3(new_n684), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n885), .A2(new_n676), .A3(new_n847), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n713), .A2(new_n444), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n846), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n630), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(G169gat), .ZN(G1348gat));
  NAND3_X1  g725(.A1(new_n924), .A2(G176gat), .A3(new_n724), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  AOI21_X1  g727(.A(G176gat), .B1(new_n924), .B2(new_n251), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n924), .A2(new_n683), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G183gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n336), .B2(new_n931), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g733(.A1(new_n924), .A2(new_n676), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(G190gat), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(G190gat), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1351gat));
  AND2_X1   g739(.A1(new_n885), .A2(new_n923), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n630), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT125), .Z(new_n944));
  AND2_X1   g743(.A1(new_n893), .A2(new_n896), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n923), .ZN(new_n946));
  OAI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n629), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n724), .A3(new_n923), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(G204gat), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(G204gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n953), .A3(new_n251), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  NAND2_X1  g754(.A1(new_n952), .A2(new_n955), .ZN(G1353gat));
  OAI21_X1  g755(.A(G211gat), .B1(new_n946), .B2(new_n655), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(KEYINPUT63), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(KEYINPUT63), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n388), .A3(new_n683), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n946), .B2(new_n684), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n389), .A3(new_n676), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


