// Benchmark "locked_c3540" written by ABC on Sat Dec 16 11:14:54 2023

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41,
    G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132,
    G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226,
    G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311,
    G317, G322, G326, G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13,
    G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124,
    G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213,
    G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283,
    G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137, new_n138, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n171, new_n172, new_n173, new_n174, new_n175,
    new_n176, new_n178, new_n179, new_n180, new_n181, new_n182, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n192, new_n193, new_n194, new_n195, new_n196, new_n197,
    new_n198, new_n199, new_n200, new_n201, new_n202, new_n203, new_n204,
    new_n205, new_n206, new_n207, new_n208, new_n209, new_n210, new_n211,
    new_n212, new_n213, new_n214, new_n215, new_n216, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223, new_n224, new_n225,
    new_n226, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978;
  NOR3_X1   g000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n137));
  INV_X1    g001(.A(G77), .ZN(new_n138));
  AND2_X1   g002(.A1(new_n137), .A2(new_n138), .ZN(G353));
  OAI21_X1  g003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g004(.A(G58), .ZN(new_n141));
  INV_X1    g005(.A(G68), .ZN(new_n142));
  NAND2_X1  g006(.A1(new_n141), .A2(new_n142), .ZN(new_n143));
  NAND2_X1  g007(.A1(new_n143), .A2(G50), .ZN(new_n144));
  INV_X1    g008(.A(G20), .ZN(new_n145));
  NAND2_X1  g009(.A1(G1), .A2(G13), .ZN(new_n146));
  NOR3_X1   g010(.A1(new_n144), .A2(new_n145), .A3(new_n146), .ZN(new_n147));
  INV_X1    g011(.A(G1), .ZN(new_n148));
  NOR2_X1   g012(.A1(new_n148), .A2(G13), .ZN(new_n149));
  NAND2_X1  g013(.A1(new_n149), .A2(G20), .ZN(new_n150));
  INV_X1    g014(.A(new_n150), .ZN(new_n151));
  OAI211_X1 g015(.A(new_n151), .B(G250), .C1(G257), .C2(G264), .ZN(new_n152));
  XNOR2_X1  g016(.A(new_n152), .B(KEYINPUT0), .ZN(new_n153));
  AOI22_X1  g017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n154));
  AOI22_X1  g018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n155));
  NAND2_X1  g019(.A1(new_n154), .A2(new_n155), .ZN(new_n156));
  AOI22_X1  g020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n157));
  AOI22_X1  g021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n158));
  NAND2_X1  g022(.A1(new_n157), .A2(new_n158), .ZN(new_n159));
  OAI22_X1  g023(.A1(new_n156), .A2(new_n159), .B1(new_n148), .B2(new_n145), .ZN(new_n160));
  OAI21_X1  g024(.A(new_n153), .B1(KEYINPUT1), .B2(new_n160), .ZN(new_n161));
  AOI211_X1 g025(.A(new_n147), .B(new_n161), .C1(KEYINPUT1), .C2(new_n160), .ZN(G361));
  XOR2_X1   g026(.A(G238), .B(G244), .Z(new_n163));
  XNOR2_X1  g027(.A(new_n163), .B(KEYINPUT2), .ZN(new_n164));
  XOR2_X1   g028(.A(G226), .B(G232), .Z(new_n165));
  XNOR2_X1  g029(.A(new_n164), .B(new_n165), .ZN(new_n166));
  XOR2_X1   g030(.A(G264), .B(G270), .Z(new_n167));
  XNOR2_X1  g031(.A(G250), .B(G257), .ZN(new_n168));
  XNOR2_X1  g032(.A(new_n167), .B(new_n168), .ZN(new_n169));
  XNOR2_X1  g033(.A(new_n166), .B(new_n169), .ZN(G358));
  XNOR2_X1  g034(.A(G50), .B(G58), .ZN(new_n171));
  XNOR2_X1  g035(.A(new_n171), .B(new_n142), .ZN(new_n172));
  XNOR2_X1  g036(.A(new_n172), .B(new_n138), .ZN(new_n173));
  XNOR2_X1  g037(.A(G87), .B(G97), .ZN(new_n174));
  XNOR2_X1  g038(.A(G107), .B(G116), .ZN(new_n175));
  XNOR2_X1  g039(.A(new_n174), .B(new_n175), .ZN(new_n176));
  XNOR2_X1  g040(.A(new_n173), .B(new_n176), .ZN(G351));
  NAND2_X1  g041(.A1(G33), .A2(G41), .ZN(new_n178));
  NAND3_X1  g042(.A1(new_n178), .A2(G1), .A3(G13), .ZN(new_n179));
  OAI21_X1  g043(.A(new_n148), .B1(G41), .B2(G45), .ZN(new_n180));
  AND2_X1   g044(.A1(new_n179), .A2(new_n180), .ZN(new_n181));
  NAND2_X1  g045(.A1(new_n181), .A2(G226), .ZN(new_n182));
  INV_X1    g046(.A(G274), .ZN(new_n183));
  NOR2_X1   g047(.A1(new_n180), .A2(new_n183), .ZN(new_n184));
  INV_X1    g048(.A(new_n184), .ZN(new_n185));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n186));
  INV_X1    g050(.A(G33), .ZN(new_n187));
  NAND2_X1  g051(.A1(new_n186), .A2(new_n187), .ZN(new_n188));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n189));
  NAND2_X1  g053(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g054(.A(G1698), .ZN(new_n191));
  NAND3_X1  g055(.A1(new_n190), .A2(G222), .A3(new_n191), .ZN(new_n192));
  NAND2_X1  g056(.A1(new_n190), .A2(G1698), .ZN(new_n193));
  INV_X1    g057(.A(G223), .ZN(new_n194));
  OAI21_X1  g058(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n196));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n197));
  NOR2_X1   g061(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g062(.A(new_n195), .B1(G77), .B2(new_n198), .ZN(new_n199));
  OAI211_X1 g063(.A(new_n182), .B(new_n185), .C1(new_n199), .C2(new_n179), .ZN(new_n200));
  NAND2_X1  g064(.A1(new_n200), .A2(G169), .ZN(new_n201));
  INV_X1    g065(.A(G179), .ZN(new_n202));
  OAI21_X1  g066(.A(new_n201), .B1(new_n202), .B2(new_n200), .ZN(new_n203));
  INV_X1    g067(.A(G13), .ZN(new_n204));
  NOR3_X1   g068(.A1(new_n204), .A2(new_n145), .A3(G1), .ZN(new_n205));
  INV_X1    g069(.A(G50), .ZN(new_n206));
  NAND2_X1  g070(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n208));
  NAND2_X1  g072(.A1(new_n208), .A2(new_n146), .ZN(new_n209));
  AOI21_X1  g073(.A(new_n209), .B1(new_n148), .B2(G20), .ZN(new_n210));
  INV_X1    g074(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g075(.A1(new_n145), .A2(new_n187), .ZN(new_n212));
  INV_X1    g076(.A(G150), .ZN(new_n213));
  OAI22_X1  g077(.A1(new_n137), .A2(new_n145), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g078(.A1(new_n187), .A2(G20), .ZN(new_n215));
  XOR2_X1   g079(.A(KEYINPUT8), .B(G58), .Z(new_n216));
  AOI21_X1  g080(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g081(.A(new_n209), .ZN(new_n218));
  OAI221_X1 g082(.A(new_n207), .B1(new_n211), .B2(new_n206), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g083(.A1(new_n203), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g084(.A1(new_n200), .A2(G200), .ZN(new_n221));
  INV_X1    g085(.A(G190), .ZN(new_n222));
  OAI21_X1  g086(.A(new_n221), .B1(new_n222), .B2(new_n200), .ZN(new_n223));
  XOR2_X1   g087(.A(new_n219), .B(KEYINPUT9), .Z(new_n224));
  OR3_X1    g088(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT10), .ZN(new_n225));
  OAI21_X1  g089(.A(KEYINPUT10), .B1(new_n223), .B2(new_n224), .ZN(new_n226));
  AOI21_X1  g090(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g091(.A(KEYINPUT7), .B1(new_n198), .B2(new_n145), .ZN(new_n228));
  NAND4_X1  g092(.A1(new_n188), .A2(KEYINPUT7), .A3(new_n145), .A4(new_n189), .ZN(new_n229));
  INV_X1    g093(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g094(.A(G68), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g095(.A(new_n212), .ZN(new_n232));
  NAND2_X1  g096(.A1(new_n232), .A2(G159), .ZN(new_n233));
  XNOR2_X1  g097(.A(G58), .B(G68), .ZN(new_n234));
  NAND2_X1  g098(.A1(new_n234), .A2(G20), .ZN(new_n235));
  NAND3_X1  g099(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g100(.A(KEYINPUT16), .ZN(new_n237));
  NAND2_X1  g101(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g102(.A1(new_n231), .A2(KEYINPUT16), .A3(new_n233), .A4(new_n235), .ZN(new_n239));
  NAND3_X1  g103(.A1(new_n238), .A2(new_n209), .A3(new_n239), .ZN(new_n240));
  INV_X1    g104(.A(new_n216), .ZN(new_n241));
  NAND2_X1  g105(.A1(new_n241), .A2(new_n205), .ZN(new_n242));
  NAND2_X1  g106(.A1(new_n210), .A2(new_n216), .ZN(new_n243));
  NAND3_X1  g107(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AND3_X1   g108(.A1(new_n179), .A2(G232), .A3(new_n180), .ZN(new_n245));
  OAI211_X1 g109(.A(G226), .B(G1698), .C1(new_n196), .C2(new_n197), .ZN(new_n246));
  OAI211_X1 g110(.A(G223), .B(new_n191), .C1(new_n196), .C2(new_n197), .ZN(new_n247));
  INV_X1    g111(.A(G87), .ZN(new_n248));
  OAI211_X1 g112(.A(new_n246), .B(new_n247), .C1(new_n187), .C2(new_n248), .ZN(new_n249));
  INV_X1    g113(.A(new_n179), .ZN(new_n250));
  AOI211_X1 g114(.A(new_n184), .B(new_n245), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g115(.A1(new_n251), .A2(G179), .ZN(new_n252));
  INV_X1    g116(.A(G169), .ZN(new_n253));
  OAI21_X1  g117(.A(new_n252), .B1(new_n253), .B2(new_n251), .ZN(new_n254));
  NAND2_X1  g118(.A1(new_n244), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g119(.A1(new_n255), .A2(KEYINPUT18), .ZN(new_n256));
  INV_X1    g120(.A(KEYINPUT18), .ZN(new_n257));
  NAND3_X1  g121(.A1(new_n244), .A2(new_n257), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g122(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g123(.A1(new_n249), .A2(new_n250), .ZN(new_n260));
  INV_X1    g124(.A(new_n245), .ZN(new_n261));
  NAND4_X1  g125(.A1(new_n260), .A2(new_n222), .A3(new_n185), .A4(new_n261), .ZN(new_n262));
  OAI21_X1  g126(.A(new_n262), .B1(new_n251), .B2(G200), .ZN(new_n263));
  NAND4_X1  g127(.A1(new_n240), .A2(new_n242), .A3(new_n263), .A4(new_n243), .ZN(new_n264));
  INV_X1    g128(.A(KEYINPUT17), .ZN(new_n265));
  XNOR2_X1  g129(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NOR2_X1   g130(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g131(.A(new_n215), .ZN(new_n268));
  NOR2_X1   g132(.A1(new_n268), .A2(new_n138), .ZN(new_n269));
  OAI22_X1  g133(.A1(new_n212), .A2(new_n206), .B1(new_n145), .B2(G68), .ZN(new_n270));
  OAI21_X1  g134(.A(new_n209), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g135(.A(new_n271), .B(KEYINPUT11), .ZN(new_n272));
  NAND2_X1  g136(.A1(new_n205), .A2(new_n142), .ZN(new_n273));
  XNOR2_X1  g137(.A(new_n273), .B(KEYINPUT12), .ZN(new_n274));
  OAI211_X1 g138(.A(new_n272), .B(new_n274), .C1(new_n142), .C2(new_n211), .ZN(new_n275));
  INV_X1    g139(.A(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g140(.A1(new_n190), .A2(G226), .A3(new_n191), .ZN(new_n277));
  NAND2_X1  g141(.A1(G33), .A2(G97), .ZN(new_n278));
  INV_X1    g142(.A(G232), .ZN(new_n279));
  OAI211_X1 g143(.A(new_n277), .B(new_n278), .C1(new_n193), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g144(.A(new_n184), .B1(new_n280), .B2(new_n250), .ZN(new_n281));
  NAND2_X1  g145(.A1(new_n181), .A2(G238), .ZN(new_n282));
  AOI21_X1  g146(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g147(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g148(.A1(new_n281), .A2(new_n276), .A3(new_n282), .ZN(new_n285));
  NAND3_X1  g149(.A1(new_n284), .A2(new_n222), .A3(new_n285), .ZN(new_n286));
  INV_X1    g150(.A(G200), .ZN(new_n287));
  AND3_X1   g151(.A1(new_n281), .A2(new_n276), .A3(new_n282), .ZN(new_n288));
  OAI21_X1  g152(.A(new_n287), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  AOI21_X1  g153(.A(new_n275), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g154(.A(G169), .B1(new_n288), .B2(new_n283), .ZN(new_n291));
  NAND2_X1  g155(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n292));
  NAND3_X1  g156(.A1(new_n284), .A2(G179), .A3(new_n285), .ZN(new_n293));
  INV_X1    g157(.A(KEYINPUT14), .ZN(new_n294));
  OAI211_X1 g158(.A(new_n294), .B(G169), .C1(new_n288), .C2(new_n283), .ZN(new_n295));
  NAND3_X1  g159(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g160(.A(new_n290), .B1(new_n296), .B2(new_n275), .ZN(new_n297));
  NAND3_X1  g161(.A1(new_n227), .A2(new_n267), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g162(.A1(new_n198), .A2(G107), .ZN(new_n299));
  INV_X1    g163(.A(G238), .ZN(new_n300));
  NAND2_X1  g164(.A1(new_n190), .A2(new_n191), .ZN(new_n301));
  OAI221_X1 g165(.A(new_n299), .B1(new_n193), .B2(new_n300), .C1(new_n279), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g166(.A1(new_n302), .A2(new_n250), .ZN(new_n303));
  AOI21_X1  g167(.A(new_n184), .B1(new_n181), .B2(G244), .ZN(new_n304));
  NAND2_X1  g168(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g169(.A1(new_n305), .A2(new_n287), .ZN(new_n306));
  OAI21_X1  g170(.A(new_n306), .B1(G190), .B2(new_n305), .ZN(new_n307));
  AOI22_X1  g171(.A1(new_n216), .A2(new_n232), .B1(G20), .B2(G77), .ZN(new_n308));
  XOR2_X1   g172(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  INV_X1    g173(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g174(.A(new_n308), .B1(new_n268), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g175(.A1(new_n311), .A2(new_n209), .B1(G77), .B2(new_n210), .ZN(new_n312));
  INV_X1    g176(.A(new_n205), .ZN(new_n313));
  OAI211_X1 g177(.A(new_n307), .B(new_n312), .C1(G77), .C2(new_n313), .ZN(new_n314));
  OAI21_X1  g178(.A(new_n312), .B1(G77), .B2(new_n313), .ZN(new_n315));
  NOR2_X1   g179(.A1(new_n305), .A2(new_n202), .ZN(new_n316));
  AOI21_X1  g180(.A(new_n253), .B1(new_n303), .B2(new_n304), .ZN(new_n317));
  OAI21_X1  g181(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g182(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g183(.A1(new_n298), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g184(.A1(new_n145), .A2(G107), .ZN(new_n321));
  XNOR2_X1  g185(.A(new_n321), .B(KEYINPUT23), .ZN(new_n322));
  NAND3_X1  g186(.A1(new_n145), .A2(G33), .A3(G116), .ZN(new_n323));
  INV_X1    g187(.A(KEYINPUT22), .ZN(new_n324));
  AOI21_X1  g188(.A(G20), .B1(new_n188), .B2(new_n189), .ZN(new_n325));
  AOI21_X1  g189(.A(new_n324), .B1(new_n325), .B2(G87), .ZN(new_n326));
  OAI211_X1 g190(.A(new_n145), .B(G87), .C1(new_n196), .C2(new_n197), .ZN(new_n327));
  NOR2_X1   g191(.A1(new_n327), .A2(KEYINPUT22), .ZN(new_n328));
  OAI211_X1 g192(.A(new_n322), .B(new_n323), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  INV_X1    g193(.A(KEYINPUT24), .ZN(new_n330));
  NAND2_X1  g194(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g195(.A(new_n327), .B(KEYINPUT22), .ZN(new_n332));
  NAND4_X1  g196(.A1(new_n332), .A2(KEYINPUT24), .A3(new_n322), .A4(new_n323), .ZN(new_n333));
  NAND3_X1  g197(.A1(new_n331), .A2(new_n333), .A3(new_n209), .ZN(new_n334));
  INV_X1    g198(.A(G107), .ZN(new_n335));
  NAND2_X1  g199(.A1(new_n205), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g200(.A(new_n336), .B(KEYINPUT25), .Z(new_n337));
  NAND2_X1  g201(.A1(new_n148), .A2(G33), .ZN(new_n338));
  NAND3_X1  g202(.A1(new_n338), .A2(new_n146), .A3(new_n208), .ZN(new_n339));
  NOR2_X1   g203(.A1(new_n339), .A2(new_n205), .ZN(new_n340));
  NAND2_X1  g204(.A1(new_n340), .A2(G107), .ZN(new_n341));
  NAND3_X1  g205(.A1(new_n334), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  OAI211_X1 g206(.A(G250), .B(new_n191), .C1(new_n196), .C2(new_n197), .ZN(new_n343));
  OAI211_X1 g207(.A(G257), .B(G1698), .C1(new_n196), .C2(new_n197), .ZN(new_n344));
  INV_X1    g208(.A(G294), .ZN(new_n345));
  OAI211_X1 g209(.A(new_n343), .B(new_n344), .C1(new_n187), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g210(.A1(new_n346), .A2(new_n250), .ZN(new_n347));
  INV_X1    g211(.A(G45), .ZN(new_n348));
  NOR2_X1   g212(.A1(new_n348), .A2(G1), .ZN(new_n349));
  NOR2_X1   g213(.A1(KEYINPUT5), .A2(G41), .ZN(new_n350));
  AND2_X1   g214(.A1(KEYINPUT5), .A2(G41), .ZN(new_n351));
  OAI211_X1 g215(.A(new_n349), .B(G274), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  OAI21_X1  g216(.A(new_n349), .B1(new_n351), .B2(new_n350), .ZN(new_n353));
  AND2_X1   g217(.A1(new_n353), .A2(new_n179), .ZN(new_n354));
  NAND2_X1  g218(.A1(new_n354), .A2(G264), .ZN(new_n355));
  NAND3_X1  g219(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g220(.A1(new_n356), .A2(G169), .ZN(new_n357));
  OAI21_X1  g221(.A(new_n357), .B1(new_n202), .B2(new_n356), .ZN(new_n358));
  NAND2_X1  g222(.A1(new_n342), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g223(.A1(new_n347), .A2(new_n355), .A3(new_n222), .A4(new_n352), .ZN(new_n360));
  AND3_X1   g224(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n361));
  OAI21_X1  g225(.A(new_n360), .B1(new_n361), .B2(G200), .ZN(new_n362));
  NAND4_X1  g226(.A1(new_n362), .A2(new_n337), .A3(new_n341), .A4(new_n334), .ZN(new_n363));
  AND2_X1   g227(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g228(.A(KEYINPUT21), .ZN(new_n365));
  OAI211_X1 g229(.A(G264), .B(G1698), .C1(new_n196), .C2(new_n197), .ZN(new_n366));
  OAI211_X1 g230(.A(G257), .B(new_n191), .C1(new_n196), .C2(new_n197), .ZN(new_n367));
  NAND3_X1  g231(.A1(new_n188), .A2(G303), .A3(new_n189), .ZN(new_n368));
  NAND3_X1  g232(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g233(.A1(new_n369), .A2(new_n250), .ZN(new_n370));
  NAND3_X1  g234(.A1(new_n353), .A2(G270), .A3(new_n179), .ZN(new_n371));
  NAND3_X1  g235(.A1(new_n370), .A2(new_n352), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g236(.A1(new_n372), .A2(G169), .ZN(new_n373));
  NOR2_X1   g237(.A1(new_n313), .A2(G116), .ZN(new_n374));
  INV_X1    g238(.A(G116), .ZN(new_n375));
  NOR3_X1   g239(.A1(new_n339), .A2(new_n205), .A3(new_n375), .ZN(new_n376));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n377));
  NOR2_X1   g241(.A1(new_n145), .A2(new_n375), .ZN(new_n378));
  NAND2_X1  g242(.A1(G33), .A2(G283), .ZN(new_n379));
  INV_X1    g243(.A(G97), .ZN(new_n380));
  OAI21_X1  g244(.A(new_n379), .B1(new_n380), .B2(G33), .ZN(new_n381));
  AOI21_X1  g245(.A(new_n378), .B1(new_n381), .B2(new_n145), .ZN(new_n382));
  OAI21_X1  g246(.A(new_n377), .B1(new_n382), .B2(new_n218), .ZN(new_n383));
  NAND2_X1  g247(.A1(new_n187), .A2(G97), .ZN(new_n384));
  AOI21_X1  g248(.A(G20), .B1(new_n384), .B2(new_n379), .ZN(new_n385));
  OAI211_X1 g249(.A(KEYINPUT20), .B(new_n209), .C1(new_n385), .C2(new_n378), .ZN(new_n386));
  AOI211_X1 g250(.A(new_n374), .B(new_n376), .C1(new_n383), .C2(new_n386), .ZN(new_n387));
  OAI21_X1  g251(.A(new_n365), .B1(new_n373), .B2(new_n387), .ZN(new_n388));
  AND4_X1   g252(.A1(new_n222), .A2(new_n370), .A3(new_n352), .A4(new_n371), .ZN(new_n389));
  INV_X1    g253(.A(new_n352), .ZN(new_n390));
  AOI21_X1  g254(.A(new_n390), .B1(new_n369), .B2(new_n250), .ZN(new_n391));
  AOI21_X1  g255(.A(G200), .B1(new_n391), .B2(new_n371), .ZN(new_n392));
  OAI21_X1  g256(.A(new_n387), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g257(.A(new_n374), .B1(new_n383), .B2(new_n386), .ZN(new_n394));
  INV_X1    g258(.A(new_n376), .ZN(new_n395));
  NAND2_X1  g259(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g260(.A1(new_n396), .A2(KEYINPUT21), .A3(G169), .A4(new_n372), .ZN(new_n397));
  INV_X1    g261(.A(new_n372), .ZN(new_n398));
  NAND3_X1  g262(.A1(new_n396), .A2(new_n398), .A3(G179), .ZN(new_n399));
  NAND4_X1  g263(.A1(new_n388), .A2(new_n393), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  OAI211_X1 g264(.A(G244), .B(new_n191), .C1(new_n196), .C2(new_n197), .ZN(new_n401));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g266(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g267(.A1(new_n190), .A2(KEYINPUT4), .A3(G244), .A4(new_n191), .ZN(new_n404));
  NAND3_X1  g268(.A1(new_n190), .A2(G250), .A3(G1698), .ZN(new_n405));
  NAND4_X1  g269(.A1(new_n403), .A2(new_n404), .A3(new_n379), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g270(.A1(new_n406), .A2(new_n250), .ZN(new_n407));
  NAND2_X1  g271(.A1(new_n354), .A2(G257), .ZN(new_n408));
  NAND3_X1  g272(.A1(new_n407), .A2(new_n352), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g273(.A1(new_n409), .A2(G169), .ZN(new_n410));
  NAND4_X1  g274(.A1(new_n407), .A2(G179), .A3(new_n352), .A4(new_n408), .ZN(new_n411));
  INV_X1    g275(.A(new_n340), .ZN(new_n412));
  NOR2_X1   g276(.A1(new_n412), .A2(new_n380), .ZN(new_n413));
  OAI21_X1  g277(.A(G107), .B1(new_n228), .B2(new_n230), .ZN(new_n414));
  NOR2_X1   g278(.A1(new_n212), .A2(new_n138), .ZN(new_n415));
  INV_X1    g279(.A(new_n415), .ZN(new_n416));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n417));
  AND2_X1   g281(.A1(G97), .A2(G107), .ZN(new_n418));
  NOR2_X1   g282(.A1(G97), .A2(G107), .ZN(new_n419));
  OAI21_X1  g283(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g284(.A1(new_n335), .A2(KEYINPUT6), .A3(G97), .ZN(new_n421));
  AOI21_X1  g285(.A(new_n145), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g286(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g287(.A1(new_n414), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g288(.A(new_n413), .B1(new_n424), .B2(new_n209), .ZN(new_n425));
  NOR2_X1   g289(.A1(new_n313), .A2(G97), .ZN(new_n426));
  INV_X1    g290(.A(new_n426), .ZN(new_n427));
  AOI22_X1  g291(.A1(new_n410), .A2(new_n411), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g292(.A(new_n413), .ZN(new_n429));
  NAND3_X1  g293(.A1(new_n188), .A2(new_n145), .A3(new_n189), .ZN(new_n430));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n431));
  NAND2_X1  g295(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g296(.A(new_n335), .B1(new_n432), .B2(new_n229), .ZN(new_n433));
  NOR3_X1   g297(.A1(new_n433), .A2(new_n415), .A3(new_n422), .ZN(new_n434));
  OAI211_X1 g298(.A(new_n427), .B(new_n429), .C1(new_n434), .C2(new_n218), .ZN(new_n435));
  NAND2_X1  g299(.A1(new_n409), .A2(new_n287), .ZN(new_n436));
  NAND4_X1  g300(.A1(new_n407), .A2(new_n222), .A3(new_n352), .A4(new_n408), .ZN(new_n437));
  AOI21_X1  g301(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g302(.A1(new_n400), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g303(.A1(new_n215), .A2(G97), .ZN(new_n440));
  XOR2_X1   g304(.A(new_n440), .B(KEYINPUT19), .Z(new_n441));
  NAND2_X1  g305(.A1(new_n325), .A2(G68), .ZN(new_n442));
  NAND2_X1  g306(.A1(new_n248), .A2(new_n380), .ZN(new_n443));
  OAI21_X1  g307(.A(G20), .B1(new_n443), .B2(G107), .ZN(new_n444));
  NAND2_X1  g308(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g309(.A(new_n209), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  OAI22_X1  g310(.A1(new_n412), .A2(new_n248), .B1(new_n313), .B2(new_n309), .ZN(new_n447));
  INV_X1    g311(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g312(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g313(.A(new_n349), .ZN(new_n450));
  NAND2_X1  g314(.A1(new_n450), .A2(G250), .ZN(new_n451));
  OAI22_X1  g315(.A1(new_n451), .A2(new_n250), .B1(new_n183), .B2(new_n450), .ZN(new_n452));
  NAND3_X1  g316(.A1(new_n190), .A2(G244), .A3(G1698), .ZN(new_n453));
  NAND2_X1  g317(.A1(G33), .A2(G116), .ZN(new_n454));
  OAI211_X1 g318(.A(new_n453), .B(new_n454), .C1(new_n301), .C2(new_n300), .ZN(new_n455));
  AOI21_X1  g319(.A(new_n452), .B1(new_n455), .B2(new_n250), .ZN(new_n456));
  NOR2_X1   g320(.A1(new_n456), .A2(new_n287), .ZN(new_n457));
  NOR2_X1   g321(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g322(.A1(new_n456), .A2(G190), .ZN(new_n459));
  NAND2_X1  g323(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g324(.A1(new_n340), .A2(new_n309), .ZN(new_n461));
  OAI211_X1 g325(.A(new_n446), .B(new_n461), .C1(new_n313), .C2(new_n309), .ZN(new_n462));
  INV_X1    g326(.A(new_n456), .ZN(new_n463));
  NAND2_X1  g327(.A1(new_n463), .A2(new_n253), .ZN(new_n464));
  NAND2_X1  g328(.A1(new_n456), .A2(new_n202), .ZN(new_n465));
  NAND3_X1  g329(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g330(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  AND4_X1   g331(.A1(new_n320), .A2(new_n364), .A3(new_n439), .A4(new_n467), .ZN(G372));
  INV_X1    g332(.A(new_n220), .ZN(new_n469));
  NAND2_X1  g333(.A1(new_n296), .A2(new_n275), .ZN(new_n470));
  INV_X1    g334(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g335(.A1(new_n227), .A2(new_n267), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g336(.A(new_n469), .B(new_n472), .C1(new_n298), .C2(new_n318), .ZN(new_n473));
  NAND2_X1  g337(.A1(new_n225), .A2(new_n226), .ZN(new_n474));
  NAND2_X1  g338(.A1(new_n474), .A2(new_n259), .ZN(new_n475));
  INV_X1    g339(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g340(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g341(.A(new_n320), .ZN(new_n478));
  INV_X1    g342(.A(new_n466), .ZN(new_n479));
  INV_X1    g343(.A(KEYINPUT26), .ZN(new_n480));
  AND3_X1   g344(.A1(new_n388), .A2(new_n397), .A3(new_n399), .ZN(new_n481));
  NAND2_X1  g345(.A1(new_n481), .A2(new_n359), .ZN(new_n482));
  AOI21_X1  g346(.A(new_n428), .B1(new_n482), .B2(new_n363), .ZN(new_n483));
  INV_X1    g347(.A(new_n460), .ZN(new_n484));
  NOR2_X1   g348(.A1(new_n484), .A2(new_n438), .ZN(new_n485));
  INV_X1    g349(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g350(.A(new_n480), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g351(.A(new_n428), .ZN(new_n488));
  NOR3_X1   g352(.A1(new_n484), .A2(new_n488), .A3(new_n480), .ZN(new_n489));
  INV_X1    g353(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g354(.A(new_n479), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g355(.A(new_n477), .B1(new_n478), .B2(new_n491), .ZN(G369));
  INV_X1    g356(.A(new_n342), .ZN(new_n493));
  NAND3_X1  g357(.A1(new_n148), .A2(new_n145), .A3(G13), .ZN(new_n494));
  OR2_X1    g358(.A1(new_n494), .A2(KEYINPUT27), .ZN(new_n495));
  NAND2_X1  g359(.A1(new_n494), .A2(KEYINPUT27), .ZN(new_n496));
  NAND3_X1  g360(.A1(new_n495), .A2(G213), .A3(new_n496), .ZN(new_n497));
  INV_X1    g361(.A(G343), .ZN(new_n498));
  NOR2_X1   g362(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g363(.A(new_n499), .ZN(new_n500));
  OAI211_X1 g364(.A(new_n359), .B(new_n363), .C1(new_n493), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g365(.A1(new_n342), .A2(new_n358), .A3(new_n499), .ZN(new_n502));
  NAND2_X1  g366(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g367(.A1(new_n481), .A2(new_n499), .ZN(new_n504));
  XNOR2_X1  g368(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g369(.A(new_n481), .ZN(new_n506));
  NOR2_X1   g370(.A1(new_n387), .A2(new_n500), .ZN(new_n507));
  NAND2_X1  g371(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g372(.A(new_n508), .B1(new_n400), .B2(new_n507), .ZN(new_n509));
  NAND2_X1  g373(.A1(new_n509), .A2(G330), .ZN(new_n510));
  NOR2_X1   g374(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g375(.A(new_n511), .ZN(new_n512));
  AOI22_X1  g376(.A1(new_n481), .A2(new_n359), .B1(new_n493), .B2(new_n362), .ZN(new_n513));
  NAND2_X1  g377(.A1(new_n513), .A2(new_n500), .ZN(new_n514));
  NAND2_X1  g378(.A1(new_n512), .A2(new_n514), .ZN(G399));
  NOR2_X1   g379(.A1(new_n150), .A2(G41), .ZN(new_n516));
  INV_X1    g380(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g381(.A1(new_n443), .A2(G107), .A3(G116), .ZN(new_n518));
  NAND3_X1  g382(.A1(new_n517), .A2(G1), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g383(.A(new_n519), .B1(new_n144), .B2(new_n517), .ZN(new_n520));
  XNOR2_X1  g384(.A(new_n520), .B(KEYINPUT28), .ZN(new_n521));
  OAI21_X1  g385(.A(KEYINPUT29), .B1(new_n491), .B2(new_n499), .ZN(new_n522));
  NAND4_X1  g386(.A1(new_n439), .A2(new_n364), .A3(new_n467), .A4(new_n500), .ZN(new_n523));
  NAND4_X1  g387(.A1(new_n456), .A2(new_n407), .A3(new_n352), .A4(new_n408), .ZN(new_n524));
  INV_X1    g388(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g389(.A1(new_n356), .A2(new_n372), .A3(new_n202), .ZN(new_n526));
  NAND3_X1  g390(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n526), .ZN(new_n527));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n528));
  NAND3_X1  g392(.A1(new_n361), .A2(new_n398), .A3(G179), .ZN(new_n529));
  OAI21_X1  g393(.A(new_n528), .B1(new_n529), .B2(new_n524), .ZN(new_n530));
  NOR2_X1   g394(.A1(new_n361), .A2(G179), .ZN(new_n531));
  NAND4_X1  g395(.A1(new_n531), .A2(new_n409), .A3(new_n372), .A4(new_n463), .ZN(new_n532));
  NAND3_X1  g396(.A1(new_n527), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g397(.A1(new_n533), .A2(KEYINPUT31), .A3(new_n499), .ZN(new_n534));
  NAND2_X1  g398(.A1(new_n533), .A2(new_n499), .ZN(new_n535));
  INV_X1    g399(.A(KEYINPUT31), .ZN(new_n536));
  NAND2_X1  g400(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g401(.A1(new_n523), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g402(.A1(new_n538), .A2(G330), .ZN(new_n539));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n540));
  OAI21_X1  g404(.A(new_n485), .B1(new_n513), .B2(new_n428), .ZN(new_n541));
  AOI21_X1  g405(.A(new_n489), .B1(new_n541), .B2(new_n480), .ZN(new_n542));
  OAI211_X1 g406(.A(new_n540), .B(new_n500), .C1(new_n542), .C2(new_n479), .ZN(new_n543));
  NAND3_X1  g407(.A1(new_n522), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  INV_X1    g408(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g409(.A(new_n521), .B1(new_n545), .B2(G1), .ZN(G364));
  NOR2_X1   g410(.A1(G13), .A2(G33), .ZN(new_n547));
  INV_X1    g411(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g412(.A1(new_n548), .A2(G20), .ZN(new_n549));
  OAI211_X1 g413(.A(new_n508), .B(new_n549), .C1(new_n400), .C2(new_n507), .ZN(new_n550));
  NOR2_X1   g414(.A1(new_n204), .A2(G20), .ZN(new_n551));
  AOI21_X1  g415(.A(new_n148), .B1(new_n551), .B2(G45), .ZN(new_n552));
  INV_X1    g416(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g417(.A1(new_n553), .A2(new_n516), .ZN(new_n554));
  NOR2_X1   g418(.A1(new_n150), .A2(new_n190), .ZN(new_n555));
  INV_X1    g419(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g420(.A(new_n556), .B1(new_n173), .B2(G45), .ZN(new_n557));
  OAI21_X1  g421(.A(new_n557), .B1(G45), .B2(new_n144), .ZN(new_n558));
  NOR2_X1   g422(.A1(new_n150), .A2(new_n198), .ZN(new_n559));
  NAND2_X1  g423(.A1(new_n559), .A2(G355), .ZN(new_n560));
  OAI211_X1 g424(.A(new_n558), .B(new_n560), .C1(G116), .C2(new_n151), .ZN(new_n561));
  AOI21_X1  g425(.A(new_n146), .B1(G20), .B2(new_n253), .ZN(new_n562));
  NOR2_X1   g426(.A1(new_n549), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g427(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NOR4_X1   g428(.A1(new_n145), .A2(new_n202), .A3(new_n222), .A4(new_n287), .ZN(new_n565));
  AOI21_X1  g429(.A(new_n190), .B1(new_n565), .B2(G326), .ZN(new_n566));
  INV_X1    g430(.A(G303), .ZN(new_n567));
  NOR2_X1   g431(.A1(new_n145), .A2(new_n287), .ZN(new_n568));
  NAND3_X1  g432(.A1(new_n568), .A2(new_n202), .A3(G190), .ZN(new_n569));
  INV_X1    g433(.A(G311), .ZN(new_n570));
  NOR4_X1   g434(.A1(new_n145), .A2(new_n202), .A3(G190), .A4(G200), .ZN(new_n571));
  INV_X1    g435(.A(new_n571), .ZN(new_n572));
  OAI221_X1 g436(.A(new_n566), .B1(new_n567), .B2(new_n569), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  NOR2_X1   g437(.A1(new_n145), .A2(new_n202), .ZN(new_n574));
  NAND3_X1  g438(.A1(new_n574), .A2(G190), .A3(new_n287), .ZN(new_n575));
  INV_X1    g439(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g440(.A1(new_n568), .A2(new_n202), .A3(new_n222), .ZN(new_n577));
  INV_X1    g441(.A(new_n577), .ZN(new_n578));
  AOI22_X1  g442(.A1(new_n576), .A2(G322), .B1(new_n578), .B2(G283), .ZN(new_n579));
  NOR2_X1   g443(.A1(G179), .A2(G200), .ZN(new_n580));
  NAND2_X1  g444(.A1(new_n580), .A2(G190), .ZN(new_n581));
  NAND2_X1  g445(.A1(new_n581), .A2(G20), .ZN(new_n582));
  INV_X1    g446(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g447(.A1(new_n574), .A2(new_n222), .A3(G200), .ZN(new_n584));
  XOR2_X1   g448(.A(KEYINPUT33), .B(G317), .Z(new_n585));
  OAI221_X1 g449(.A(new_n579), .B1(new_n345), .B2(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g450(.A1(new_n580), .A2(G20), .A3(new_n222), .ZN(new_n587));
  INV_X1    g451(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g452(.A(new_n573), .B(new_n586), .C1(G329), .C2(new_n588), .ZN(new_n589));
  INV_X1    g453(.A(new_n569), .ZN(new_n590));
  NAND2_X1  g454(.A1(new_n590), .A2(G87), .ZN(new_n591));
  OAI221_X1 g455(.A(new_n591), .B1(new_n141), .B2(new_n575), .C1(new_n335), .C2(new_n577), .ZN(new_n592));
  INV_X1    g456(.A(new_n584), .ZN(new_n593));
  AOI22_X1  g457(.A1(new_n593), .A2(G68), .B1(new_n565), .B2(G50), .ZN(new_n594));
  OAI21_X1  g458(.A(new_n594), .B1(new_n380), .B2(new_n583), .ZN(new_n595));
  NAND2_X1  g459(.A1(new_n588), .A2(G159), .ZN(new_n596));
  XNOR2_X1  g460(.A(new_n596), .B(KEYINPUT32), .ZN(new_n597));
  OAI21_X1  g461(.A(new_n190), .B1(new_n572), .B2(new_n138), .ZN(new_n598));
  NOR4_X1   g462(.A1(new_n592), .A2(new_n595), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  OAI21_X1  g463(.A(new_n562), .B1(new_n589), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g464(.A1(new_n550), .A2(new_n554), .A3(new_n564), .A4(new_n600), .ZN(new_n601));
  INV_X1    g465(.A(new_n554), .ZN(new_n602));
  NAND2_X1  g466(.A1(new_n510), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g467(.A1(new_n509), .A2(G330), .ZN(new_n604));
  OAI21_X1  g468(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(G396));
  NAND2_X1  g469(.A1(new_n578), .A2(G68), .ZN(new_n606));
  OAI221_X1 g470(.A(new_n606), .B1(new_n206), .B2(new_n569), .C1(new_n141), .C2(new_n583), .ZN(new_n607));
  INV_X1    g471(.A(G132), .ZN(new_n608));
  AOI22_X1  g472(.A1(new_n576), .A2(G143), .B1(new_n571), .B2(G159), .ZN(new_n609));
  INV_X1    g473(.A(G137), .ZN(new_n610));
  INV_X1    g474(.A(new_n565), .ZN(new_n611));
  OAI221_X1 g475(.A(new_n609), .B1(new_n610), .B2(new_n611), .C1(new_n213), .C2(new_n584), .ZN(new_n612));
  INV_X1    g476(.A(KEYINPUT34), .ZN(new_n613));
  OAI221_X1 g477(.A(new_n190), .B1(new_n608), .B2(new_n587), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  AOI211_X1 g478(.A(new_n607), .B(new_n614), .C1(new_n613), .C2(new_n612), .ZN(new_n615));
  AOI22_X1  g479(.A1(G97), .A2(new_n582), .B1(new_n571), .B2(G116), .ZN(new_n616));
  INV_X1    g480(.A(G283), .ZN(new_n617));
  OAI221_X1 g481(.A(new_n616), .B1(new_n617), .B2(new_n584), .C1(new_n345), .C2(new_n575), .ZN(new_n618));
  OAI21_X1  g482(.A(new_n198), .B1(new_n611), .B2(new_n567), .ZN(new_n619));
  NOR2_X1   g483(.A1(new_n587), .A2(new_n570), .ZN(new_n620));
  OAI22_X1  g484(.A1(new_n577), .A2(new_n248), .B1(new_n569), .B2(new_n335), .ZN(new_n621));
  NOR4_X1   g485(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  OAI21_X1  g486(.A(new_n562), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g487(.A1(new_n562), .A2(new_n547), .ZN(new_n624));
  AOI21_X1  g488(.A(new_n602), .B1(new_n138), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g489(.A1(new_n318), .A2(new_n315), .A3(new_n499), .ZN(new_n626));
  NAND2_X1  g490(.A1(new_n315), .A2(new_n499), .ZN(new_n627));
  AOI21_X1  g491(.A(new_n626), .B1(new_n319), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g492(.A(new_n623), .B(new_n625), .C1(new_n628), .C2(new_n548), .ZN(new_n629));
  INV_X1    g493(.A(new_n319), .ZN(new_n630));
  OAI211_X1 g494(.A(new_n630), .B(new_n500), .C1(new_n542), .C2(new_n479), .ZN(new_n631));
  NOR2_X1   g495(.A1(new_n491), .A2(new_n499), .ZN(new_n632));
  OAI21_X1  g496(.A(new_n631), .B1(new_n632), .B2(new_n628), .ZN(new_n633));
  XNOR2_X1  g497(.A(new_n633), .B(new_n539), .ZN(new_n634));
  OAI21_X1  g498(.A(new_n629), .B1(new_n634), .B2(new_n554), .ZN(G384));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n636));
  INV_X1    g500(.A(new_n497), .ZN(new_n637));
  NAND2_X1  g501(.A1(new_n244), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g502(.A1(new_n244), .A2(new_n257), .A3(new_n254), .ZN(new_n639));
  AOI21_X1  g503(.A(new_n257), .B1(new_n244), .B2(new_n254), .ZN(new_n640));
  NOR2_X1   g504(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g505(.A(new_n264), .B(KEYINPUT17), .ZN(new_n642));
  AOI21_X1  g506(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g507(.A(new_n244), .B1(new_n254), .B2(new_n637), .ZN(new_n644));
  INV_X1    g508(.A(KEYINPUT37), .ZN(new_n645));
  AND3_X1   g509(.A1(new_n644), .A2(new_n645), .A3(new_n264), .ZN(new_n646));
  AOI21_X1  g510(.A(new_n645), .B1(new_n644), .B2(new_n264), .ZN(new_n647));
  NOR2_X1   g511(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g512(.A(new_n636), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  INV_X1    g513(.A(new_n638), .ZN(new_n650));
  OAI21_X1  g514(.A(new_n650), .B1(new_n259), .B2(new_n266), .ZN(new_n651));
  NAND2_X1  g515(.A1(new_n644), .A2(new_n264), .ZN(new_n652));
  NAND2_X1  g516(.A1(new_n652), .A2(KEYINPUT37), .ZN(new_n653));
  NAND3_X1  g517(.A1(new_n644), .A2(new_n645), .A3(new_n264), .ZN(new_n654));
  NAND2_X1  g518(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g519(.A1(new_n651), .A2(new_n655), .A3(KEYINPUT38), .ZN(new_n656));
  NAND2_X1  g520(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  INV_X1    g521(.A(new_n290), .ZN(new_n658));
  NAND2_X1  g522(.A1(new_n275), .A2(new_n499), .ZN(new_n659));
  NAND3_X1  g523(.A1(new_n470), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g524(.A(new_n660), .B1(new_n470), .B2(new_n500), .ZN(new_n661));
  AND2_X1   g525(.A1(new_n538), .A2(new_n628), .ZN(new_n662));
  AND4_X1   g526(.A1(KEYINPUT40), .A2(new_n657), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  AOI22_X1  g527(.A1(new_n471), .A2(new_n499), .B1(new_n297), .B2(new_n659), .ZN(new_n664));
  AOI21_X1  g528(.A(new_n664), .B1(new_n649), .B2(new_n656), .ZN(new_n665));
  AOI21_X1  g529(.A(KEYINPUT40), .B1(new_n665), .B2(new_n662), .ZN(new_n666));
  NOR2_X1   g530(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g531(.A1(new_n320), .A2(new_n538), .ZN(new_n668));
  XNOR2_X1  g532(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g533(.A1(new_n669), .A2(G330), .ZN(new_n670));
  AOI21_X1  g534(.A(new_n478), .B1(new_n522), .B2(new_n543), .ZN(new_n671));
  NOR3_X1   g535(.A1(new_n671), .A2(new_n476), .A3(new_n473), .ZN(new_n672));
  NOR2_X1   g536(.A1(new_n641), .A2(new_n637), .ZN(new_n673));
  OR2_X1    g537(.A1(new_n318), .A2(new_n499), .ZN(new_n674));
  NAND2_X1  g538(.A1(new_n631), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g539(.A(new_n673), .B1(new_n675), .B2(new_n665), .ZN(new_n676));
  INV_X1    g540(.A(KEYINPUT39), .ZN(new_n677));
  NOR3_X1   g541(.A1(new_n643), .A2(new_n648), .A3(new_n636), .ZN(new_n678));
  AOI21_X1  g542(.A(KEYINPUT38), .B1(new_n651), .B2(new_n655), .ZN(new_n679));
  OAI21_X1  g543(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g544(.A1(new_n649), .A2(KEYINPUT39), .A3(new_n656), .ZN(new_n681));
  NAND4_X1  g545(.A1(new_n680), .A2(new_n471), .A3(new_n500), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g546(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g547(.A(new_n672), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g548(.A(new_n670), .B(new_n684), .ZN(new_n685));
  OAI21_X1  g549(.A(new_n685), .B1(new_n148), .B2(new_n551), .ZN(new_n686));
  NAND2_X1  g550(.A1(new_n420), .A2(new_n421), .ZN(new_n687));
  AOI21_X1  g551(.A(new_n375), .B1(new_n687), .B2(KEYINPUT35), .ZN(new_n688));
  NOR2_X1   g552(.A1(new_n146), .A2(new_n145), .ZN(new_n689));
  OAI211_X1 g553(.A(new_n688), .B(new_n689), .C1(KEYINPUT35), .C2(new_n687), .ZN(new_n690));
  XNOR2_X1  g554(.A(new_n690), .B(KEYINPUT36), .ZN(new_n691));
  NAND2_X1  g555(.A1(new_n172), .A2(G77), .ZN(new_n692));
  NAND2_X1  g556(.A1(new_n692), .A2(G50), .ZN(new_n693));
  OAI211_X1 g557(.A(new_n693), .B(new_n149), .C1(G50), .C2(G68), .ZN(new_n694));
  NAND3_X1  g558(.A1(new_n686), .A2(new_n691), .A3(new_n694), .ZN(G367));
  NOR2_X1   g559(.A1(new_n569), .A2(new_n141), .ZN(new_n696));
  NAND2_X1  g560(.A1(new_n565), .A2(G143), .ZN(new_n697));
  NAND2_X1  g561(.A1(new_n582), .A2(G68), .ZN(new_n698));
  OAI211_X1 g562(.A(new_n697), .B(new_n698), .C1(new_n213), .C2(new_n575), .ZN(new_n699));
  AOI211_X1 g563(.A(new_n696), .B(new_n699), .C1(G137), .C2(new_n588), .ZN(new_n700));
  NAND2_X1  g564(.A1(new_n593), .A2(G159), .ZN(new_n701));
  NAND2_X1  g565(.A1(new_n578), .A2(G77), .ZN(new_n702));
  AOI21_X1  g566(.A(new_n198), .B1(new_n571), .B2(G50), .ZN(new_n703));
  NAND4_X1  g567(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g568(.A1(new_n577), .A2(new_n380), .ZN(new_n705));
  OR3_X1    g569(.A1(new_n569), .A2(KEYINPUT46), .A3(new_n375), .ZN(new_n706));
  OAI21_X1  g570(.A(KEYINPUT46), .B1(new_n569), .B2(new_n375), .ZN(new_n707));
  AOI21_X1  g571(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g572(.A(new_n708), .B1(new_n570), .B2(new_n611), .ZN(new_n709));
  AOI21_X1  g573(.A(new_n709), .B1(G283), .B2(new_n571), .ZN(new_n710));
  OAI221_X1 g574(.A(new_n710), .B1(new_n335), .B2(new_n583), .C1(new_n567), .C2(new_n575), .ZN(new_n711));
  INV_X1    g575(.A(G317), .ZN(new_n712));
  OAI221_X1 g576(.A(new_n198), .B1(new_n587), .B2(new_n712), .C1(new_n584), .C2(new_n345), .ZN(new_n713));
  OAI21_X1  g577(.A(new_n704), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g578(.A(new_n714), .B(KEYINPUT47), .ZN(new_n715));
  NAND2_X1  g579(.A1(new_n715), .A2(new_n562), .ZN(new_n716));
  NAND2_X1  g580(.A1(new_n449), .A2(new_n499), .ZN(new_n717));
  NOR2_X1   g581(.A1(new_n466), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g582(.A(new_n718), .B1(new_n467), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g583(.A1(new_n719), .A2(new_n549), .ZN(new_n720));
  OAI221_X1 g584(.A(new_n563), .B1(new_n151), .B2(new_n310), .C1(new_n169), .C2(new_n556), .ZN(new_n721));
  NAND4_X1  g585(.A1(new_n716), .A2(new_n554), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  INV_X1    g586(.A(new_n438), .ZN(new_n723));
  NAND2_X1  g587(.A1(new_n435), .A2(new_n499), .ZN(new_n724));
  NAND3_X1  g588(.A1(new_n488), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g589(.A1(new_n428), .A2(new_n499), .ZN(new_n726));
  NAND2_X1  g590(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g591(.A1(new_n727), .A2(new_n503), .A3(new_n504), .ZN(new_n728));
  OR2_X1    g592(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n729));
  OAI21_X1  g593(.A(new_n488), .B1(new_n359), .B2(new_n438), .ZN(new_n730));
  NAND2_X1  g594(.A1(new_n730), .A2(new_n500), .ZN(new_n731));
  NAND2_X1  g595(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n732));
  NAND3_X1  g596(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g597(.A(KEYINPUT43), .ZN(new_n734));
  NAND2_X1  g598(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g599(.A1(new_n511), .A2(new_n727), .ZN(new_n736));
  XNOR2_X1  g600(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g601(.A(new_n719), .B1(new_n733), .B2(new_n734), .ZN(new_n738));
  XOR2_X1   g602(.A(new_n737), .B(new_n738), .Z(new_n739));
  NOR2_X1   g603(.A1(new_n514), .A2(new_n727), .ZN(new_n740));
  XNOR2_X1  g604(.A(new_n740), .B(KEYINPUT44), .ZN(new_n741));
  AND2_X1   g605(.A1(new_n514), .A2(new_n727), .ZN(new_n742));
  NOR2_X1   g606(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n743));
  AND2_X1   g607(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n744));
  OAI21_X1  g608(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g609(.A1(new_n745), .A2(new_n511), .ZN(new_n746));
  OAI211_X1 g610(.A(new_n512), .B(new_n741), .C1(new_n743), .C2(new_n744), .ZN(new_n747));
  NAND2_X1  g611(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g612(.A(new_n505), .B(new_n510), .ZN(new_n749));
  OAI21_X1  g613(.A(new_n545), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g614(.A(new_n516), .B(KEYINPUT41), .ZN(new_n751));
  AOI21_X1  g615(.A(new_n553), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g616(.A(new_n722), .B1(new_n739), .B2(new_n752), .ZN(G387));
  OR2_X1    g617(.A1(new_n544), .A2(new_n749), .ZN(new_n754));
  AOI21_X1  g618(.A(new_n517), .B1(new_n544), .B2(new_n749), .ZN(new_n755));
  NAND2_X1  g619(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g620(.A(new_n198), .B1(new_n577), .B2(new_n375), .ZN(new_n757));
  AOI22_X1  g621(.A1(new_n565), .A2(G322), .B1(new_n571), .B2(G303), .ZN(new_n758));
  OAI221_X1 g622(.A(new_n758), .B1(new_n570), .B2(new_n584), .C1(new_n712), .C2(new_n575), .ZN(new_n759));
  INV_X1    g623(.A(KEYINPUT48), .ZN(new_n760));
  AOI22_X1  g624(.A1(new_n759), .A2(new_n760), .B1(G294), .B2(new_n590), .ZN(new_n761));
  OAI221_X1 g625(.A(new_n761), .B1(new_n760), .B2(new_n759), .C1(new_n617), .C2(new_n583), .ZN(new_n762));
  XOR2_X1   g626(.A(new_n762), .B(KEYINPUT49), .Z(new_n763));
  AOI211_X1 g627(.A(new_n757), .B(new_n763), .C1(G326), .C2(new_n588), .ZN(new_n764));
  NAND2_X1  g628(.A1(new_n590), .A2(G77), .ZN(new_n765));
  INV_X1    g629(.A(G159), .ZN(new_n766));
  OAI221_X1 g630(.A(new_n765), .B1(new_n206), .B2(new_n575), .C1(new_n766), .C2(new_n611), .ZN(new_n767));
  AOI21_X1  g631(.A(new_n767), .B1(G150), .B2(new_n588), .ZN(new_n768));
  OAI221_X1 g632(.A(new_n768), .B1(new_n142), .B2(new_n572), .C1(new_n310), .C2(new_n583), .ZN(new_n769));
  NOR2_X1   g633(.A1(new_n241), .A2(new_n584), .ZN(new_n770));
  NOR4_X1   g634(.A1(new_n769), .A2(new_n198), .A3(new_n705), .A4(new_n770), .ZN(new_n771));
  OAI21_X1  g635(.A(new_n562), .B1(new_n764), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g636(.A1(new_n166), .A2(new_n348), .ZN(new_n773));
  INV_X1    g637(.A(new_n518), .ZN(new_n774));
  AOI22_X1  g638(.A1(new_n773), .A2(new_n555), .B1(new_n774), .B2(new_n559), .ZN(new_n775));
  NAND2_X1  g639(.A1(new_n216), .A2(new_n206), .ZN(new_n776));
  OAI221_X1 g640(.A(new_n518), .B1(new_n142), .B2(new_n138), .C1(new_n776), .C2(KEYINPUT50), .ZN(new_n777));
  AOI211_X1 g641(.A(G45), .B(new_n777), .C1(KEYINPUT50), .C2(new_n776), .ZN(new_n778));
  OAI22_X1  g642(.A1(new_n775), .A2(new_n778), .B1(G107), .B2(new_n151), .ZN(new_n779));
  NAND2_X1  g643(.A1(new_n779), .A2(new_n563), .ZN(new_n780));
  NAND3_X1  g644(.A1(new_n501), .A2(new_n502), .A3(new_n549), .ZN(new_n781));
  NAND4_X1  g645(.A1(new_n772), .A2(new_n554), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  OAI211_X1 g646(.A(new_n756), .B(new_n782), .C1(new_n552), .C2(new_n749), .ZN(G393));
  OR2_X1    g647(.A1(new_n754), .A2(new_n748), .ZN(new_n784));
  AOI21_X1  g648(.A(new_n517), .B1(new_n754), .B2(new_n748), .ZN(new_n785));
  AND2_X1   g649(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g650(.A1(new_n611), .A2(new_n213), .B1(new_n766), .B2(new_n575), .ZN(new_n787));
  XNOR2_X1  g651(.A(new_n787), .B(KEYINPUT51), .ZN(new_n788));
  OAI221_X1 g652(.A(new_n788), .B1(new_n142), .B2(new_n569), .C1(new_n241), .C2(new_n572), .ZN(new_n789));
  AOI22_X1  g653(.A1(G50), .A2(new_n593), .B1(new_n578), .B2(G87), .ZN(new_n790));
  AOI21_X1  g654(.A(new_n198), .B1(new_n588), .B2(G143), .ZN(new_n791));
  OAI211_X1 g655(.A(new_n790), .B(new_n791), .C1(new_n138), .C2(new_n583), .ZN(new_n792));
  OAI22_X1  g656(.A1(new_n611), .A2(new_n712), .B1(new_n570), .B2(new_n575), .ZN(new_n793));
  XNOR2_X1  g657(.A(new_n793), .B(KEYINPUT52), .ZN(new_n794));
  OAI21_X1  g658(.A(new_n794), .B1(new_n375), .B2(new_n583), .ZN(new_n795));
  NOR2_X1   g659(.A1(new_n584), .A2(new_n567), .ZN(new_n796));
  OAI21_X1  g660(.A(new_n198), .B1(new_n577), .B2(new_n335), .ZN(new_n797));
  AOI211_X1 g661(.A(new_n796), .B(new_n797), .C1(G322), .C2(new_n588), .ZN(new_n798));
  OAI221_X1 g662(.A(new_n798), .B1(new_n617), .B2(new_n569), .C1(new_n345), .C2(new_n572), .ZN(new_n799));
  OAI22_X1  g663(.A1(new_n789), .A2(new_n792), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g664(.A1(new_n800), .A2(new_n562), .ZN(new_n801));
  NAND2_X1  g665(.A1(new_n176), .A2(new_n555), .ZN(new_n802));
  AOI211_X1 g666(.A(new_n562), .B(new_n549), .C1(G97), .C2(new_n150), .ZN(new_n803));
  AOI21_X1  g667(.A(new_n602), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g668(.A(new_n549), .ZN(new_n805));
  OAI211_X1 g669(.A(new_n801), .B(new_n804), .C1(new_n727), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g670(.A(new_n806), .B1(new_n748), .B2(new_n552), .ZN(new_n807));
  OR2_X1    g671(.A1(new_n786), .A2(new_n807), .ZN(G390));
  OAI21_X1  g672(.A(new_n628), .B1(new_n542), .B2(new_n479), .ZN(new_n809));
  NAND3_X1  g673(.A1(new_n809), .A2(new_n470), .A3(new_n318), .ZN(new_n810));
  NOR2_X1   g674(.A1(new_n290), .A2(new_n499), .ZN(new_n811));
  NAND4_X1  g675(.A1(new_n810), .A2(new_n680), .A3(new_n681), .A4(new_n811), .ZN(new_n812));
  INV_X1    g676(.A(new_n812), .ZN(new_n813));
  NAND4_X1  g677(.A1(new_n661), .A2(G330), .A3(new_n538), .A4(new_n628), .ZN(new_n814));
  INV_X1    g678(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g679(.A(new_n657), .B1(new_n810), .B2(new_n811), .ZN(new_n816));
  NOR3_X1   g680(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g681(.A(new_n816), .ZN(new_n818));
  AOI21_X1  g682(.A(new_n814), .B1(new_n818), .B2(new_n812), .ZN(new_n819));
  NOR2_X1   g683(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g684(.A1(new_n544), .A2(new_n320), .ZN(new_n821));
  NAND3_X1  g685(.A1(new_n538), .A2(G330), .A3(new_n628), .ZN(new_n822));
  NAND2_X1  g686(.A1(new_n822), .A2(new_n664), .ZN(new_n823));
  NAND2_X1  g687(.A1(new_n823), .A2(new_n814), .ZN(new_n824));
  NAND3_X1  g688(.A1(new_n824), .A2(new_n631), .A3(new_n674), .ZN(new_n825));
  NAND3_X1  g689(.A1(new_n675), .A2(new_n814), .A3(new_n823), .ZN(new_n826));
  NAND4_X1  g690(.A1(new_n821), .A2(new_n477), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g691(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g692(.A(new_n820), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g693(.A1(new_n829), .A2(new_n516), .ZN(new_n830));
  NAND2_X1  g694(.A1(new_n680), .A2(new_n681), .ZN(new_n831));
  NAND2_X1  g695(.A1(new_n831), .A2(new_n547), .ZN(new_n832));
  NOR2_X1   g696(.A1(new_n569), .A2(new_n213), .ZN(new_n833));
  OR2_X1    g697(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n834));
  NAND2_X1  g698(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g699(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g700(.A(new_n836), .B1(new_n206), .B2(new_n577), .ZN(new_n837));
  AOI21_X1  g701(.A(new_n837), .B1(G128), .B2(new_n565), .ZN(new_n838));
  NAND2_X1  g702(.A1(new_n588), .A2(G125), .ZN(new_n839));
  XOR2_X1   g703(.A(KEYINPUT54), .B(G143), .Z(new_n840));
  INV_X1    g704(.A(new_n840), .ZN(new_n841));
  OAI221_X1 g705(.A(new_n839), .B1(new_n608), .B2(new_n575), .C1(new_n572), .C2(new_n841), .ZN(new_n842));
  AOI211_X1 g706(.A(new_n198), .B(new_n842), .C1(G137), .C2(new_n593), .ZN(new_n843));
  OAI211_X1 g707(.A(new_n838), .B(new_n843), .C1(new_n766), .C2(new_n583), .ZN(new_n844));
  INV_X1    g708(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g709(.A1(new_n576), .A2(G116), .ZN(new_n846));
  NAND2_X1  g710(.A1(new_n565), .A2(G283), .ZN(new_n847));
  NAND4_X1  g711(.A1(new_n591), .A2(new_n606), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI22_X1  g712(.A1(G294), .A2(new_n588), .B1(new_n571), .B2(G97), .ZN(new_n849));
  OAI21_X1  g713(.A(new_n849), .B1(new_n335), .B2(new_n584), .ZN(new_n850));
  NOR2_X1   g714(.A1(new_n583), .A2(new_n138), .ZN(new_n851));
  NOR4_X1   g715(.A1(new_n848), .A2(new_n850), .A3(new_n190), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g716(.A(new_n562), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g717(.A(new_n602), .B1(new_n241), .B2(new_n624), .ZN(new_n854));
  NAND3_X1  g718(.A1(new_n832), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g719(.A(new_n855), .B1(new_n820), .B2(new_n552), .ZN(new_n856));
  INV_X1    g720(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g721(.A1(new_n830), .A2(new_n857), .ZN(G378));
  NAND3_X1  g722(.A1(new_n683), .A2(new_n667), .A3(G330), .ZN(new_n859));
  OAI211_X1 g723(.A(new_n662), .B(new_n661), .C1(new_n678), .C2(new_n679), .ZN(new_n860));
  INV_X1    g724(.A(KEYINPUT40), .ZN(new_n861));
  NAND2_X1  g725(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g726(.A1(new_n665), .A2(KEYINPUT40), .A3(new_n662), .ZN(new_n863));
  NAND3_X1  g727(.A1(new_n862), .A2(G330), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g728(.A1(new_n864), .A2(new_n676), .A3(new_n682), .ZN(new_n865));
  NAND2_X1  g729(.A1(new_n219), .A2(new_n637), .ZN(new_n866));
  XNOR2_X1  g730(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  XNOR2_X1  g731(.A(new_n867), .B(KEYINPUT56), .ZN(new_n868));
  XNOR2_X1  g732(.A(new_n227), .B(new_n868), .ZN(new_n869));
  AND3_X1   g733(.A1(new_n859), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g734(.A(new_n869), .B1(new_n859), .B2(new_n865), .ZN(new_n871));
  OAI21_X1  g735(.A(new_n815), .B1(new_n813), .B2(new_n816), .ZN(new_n872));
  NAND3_X1  g736(.A1(new_n818), .A2(new_n814), .A3(new_n812), .ZN(new_n873));
  AOI21_X1  g737(.A(new_n827), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g738(.A1(new_n821), .A2(new_n477), .ZN(new_n875));
  OAI22_X1  g739(.A1(new_n870), .A2(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g740(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n877));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n878));
  OAI221_X1 g742(.A(new_n878), .B1(new_n874), .B2(new_n875), .C1(new_n870), .C2(new_n871), .ZN(new_n879));
  NAND2_X1  g743(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g744(.A1(new_n880), .A2(new_n516), .ZN(new_n881));
  NAND2_X1  g745(.A1(new_n869), .A2(new_n547), .ZN(new_n882));
  NOR2_X1   g746(.A1(new_n575), .A2(new_n335), .ZN(new_n883));
  AOI22_X1  g747(.A1(new_n578), .A2(G58), .B1(new_n309), .B2(new_n571), .ZN(new_n884));
  OAI221_X1 g748(.A(new_n884), .B1(new_n375), .B2(new_n611), .C1(new_n617), .C2(new_n587), .ZN(new_n885));
  AOI211_X1 g749(.A(new_n883), .B(new_n885), .C1(G97), .C2(new_n593), .ZN(new_n886));
  NOR2_X1   g750(.A1(new_n190), .A2(G41), .ZN(new_n887));
  NAND4_X1  g751(.A1(new_n886), .A2(new_n698), .A3(new_n765), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g752(.A(new_n888), .B(KEYINPUT58), .Z(new_n889));
  OAI22_X1  g753(.A1(new_n841), .A2(new_n569), .B1(new_n608), .B2(new_n584), .ZN(new_n890));
  AOI22_X1  g754(.A1(G150), .A2(new_n582), .B1(new_n571), .B2(G137), .ZN(new_n891));
  INV_X1    g755(.A(G128), .ZN(new_n892));
  OAI21_X1  g756(.A(new_n891), .B1(new_n892), .B2(new_n575), .ZN(new_n893));
  AOI211_X1 g757(.A(new_n890), .B(new_n893), .C1(G125), .C2(new_n565), .ZN(new_n894));
  XNOR2_X1  g758(.A(new_n894), .B(KEYINPUT59), .ZN(new_n895));
  AOI211_X1 g759(.A(G33), .B(G41), .C1(new_n588), .C2(G124), .ZN(new_n896));
  OAI211_X1 g760(.A(new_n895), .B(new_n896), .C1(new_n766), .C2(new_n577), .ZN(new_n897));
  OAI21_X1  g761(.A(new_n206), .B1(G33), .B2(G41), .ZN(new_n898));
  OAI21_X1  g762(.A(new_n897), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g763(.A(new_n562), .B1(new_n889), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g764(.A1(new_n624), .A2(new_n206), .ZN(new_n901));
  NAND4_X1  g765(.A1(new_n882), .A2(new_n554), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g766(.A(new_n902), .ZN(new_n903));
  OR2_X1    g767(.A1(new_n870), .A2(new_n871), .ZN(new_n904));
  AOI21_X1  g768(.A(new_n903), .B1(new_n904), .B2(new_n553), .ZN(new_n905));
  NAND2_X1  g769(.A1(new_n881), .A2(new_n905), .ZN(G375));
  NAND2_X1  g770(.A1(new_n825), .A2(new_n826), .ZN(new_n907));
  NAND2_X1  g771(.A1(new_n875), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g772(.A1(new_n908), .A2(new_n751), .A3(new_n827), .ZN(new_n909));
  NAND3_X1  g773(.A1(new_n825), .A2(new_n553), .A3(new_n826), .ZN(new_n910));
  AOI22_X1  g774(.A1(G303), .A2(new_n588), .B1(new_n571), .B2(G107), .ZN(new_n911));
  OAI211_X1 g775(.A(new_n911), .B(new_n198), .C1(new_n345), .C2(new_n611), .ZN(new_n912));
  AOI22_X1  g776(.A1(G97), .A2(new_n590), .B1(new_n593), .B2(G116), .ZN(new_n913));
  OAI211_X1 g777(.A(new_n913), .B(new_n702), .C1(new_n617), .C2(new_n575), .ZN(new_n914));
  AOI211_X1 g778(.A(new_n912), .B(new_n914), .C1(new_n309), .C2(new_n582), .ZN(new_n915));
  AOI22_X1  g779(.A1(new_n593), .A2(new_n840), .B1(G150), .B2(new_n571), .ZN(new_n916));
  OAI221_X1 g780(.A(new_n916), .B1(new_n141), .B2(new_n577), .C1(new_n610), .C2(new_n575), .ZN(new_n917));
  NOR2_X1   g781(.A1(new_n583), .A2(new_n206), .ZN(new_n918));
  NOR2_X1   g782(.A1(new_n569), .A2(new_n766), .ZN(new_n919));
  OAI221_X1 g783(.A(new_n190), .B1(new_n587), .B2(new_n892), .C1(new_n611), .C2(new_n608), .ZN(new_n920));
  NOR4_X1   g784(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g785(.A(new_n562), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g786(.A(new_n602), .B1(new_n142), .B2(new_n624), .ZN(new_n923));
  OAI211_X1 g787(.A(new_n922), .B(new_n923), .C1(new_n661), .C2(new_n548), .ZN(new_n924));
  AND2_X1   g788(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g789(.A1(new_n909), .A2(new_n925), .ZN(G381));
  AOI21_X1  g790(.A(new_n856), .B1(new_n829), .B2(new_n516), .ZN(new_n927));
  NAND3_X1  g791(.A1(new_n881), .A2(new_n927), .A3(new_n905), .ZN(new_n928));
  INV_X1    g792(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g793(.A1(G381), .A2(G384), .ZN(new_n930));
  NOR2_X1   g794(.A1(new_n786), .A2(new_n807), .ZN(new_n931));
  OAI211_X1 g795(.A(new_n931), .B(new_n722), .C1(new_n739), .C2(new_n752), .ZN(new_n932));
  NOR3_X1   g796(.A1(new_n932), .A2(G396), .A3(G393), .ZN(new_n933));
  NAND3_X1  g797(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(G407));
  OAI211_X1 g798(.A(G407), .B(G213), .C1(G343), .C2(new_n928), .ZN(G409));
  AND2_X1   g799(.A1(new_n908), .A2(KEYINPUT60), .ZN(new_n936));
  NOR2_X1   g800(.A1(new_n908), .A2(KEYINPUT60), .ZN(new_n937));
  OAI211_X1 g801(.A(new_n516), .B(new_n827), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  AND3_X1   g802(.A1(new_n938), .A2(G384), .A3(new_n925), .ZN(new_n939));
  AOI21_X1  g803(.A(G384), .B1(new_n938), .B2(new_n925), .ZN(new_n940));
  OR2_X1    g804(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g805(.A1(new_n498), .A2(G213), .A3(G2897), .ZN(new_n942));
  NOR2_X1   g806(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g807(.A1(G390), .A2(G387), .ZN(new_n944));
  XOR2_X1   g808(.A(G393), .B(G396), .Z(new_n945));
  AND3_X1   g809(.A1(new_n932), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g810(.A(new_n945), .B1(new_n932), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g811(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g812(.A(new_n517), .B1(new_n877), .B2(new_n879), .ZN(new_n949));
  NAND2_X1  g813(.A1(new_n904), .A2(new_n553), .ZN(new_n950));
  NAND2_X1  g814(.A1(new_n950), .A2(new_n902), .ZN(new_n951));
  OAI21_X1  g815(.A(G378), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g816(.A1(new_n498), .A2(G213), .ZN(new_n953));
  INV_X1    g817(.A(new_n751), .ZN(new_n954));
  OAI211_X1 g818(.A(new_n927), .B(new_n905), .C1(new_n954), .C2(new_n876), .ZN(new_n955));
  NOR2_X1   g819(.A1(new_n939), .A2(new_n940), .ZN(new_n956));
  NAND4_X1  g820(.A1(new_n952), .A2(new_n953), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  INV_X1    g821(.A(KEYINPUT63), .ZN(new_n958));
  AOI211_X1 g822(.A(new_n943), .B(new_n948), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND4_X1   g823(.A1(new_n953), .A2(new_n952), .A3(new_n955), .A4(new_n956), .ZN(new_n960));
  AOI21_X1  g824(.A(KEYINPUT61), .B1(new_n960), .B2(KEYINPUT63), .ZN(new_n961));
  NAND3_X1  g825(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n962));
  INV_X1    g826(.A(new_n942), .ZN(new_n963));
  NOR2_X1   g827(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g828(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g829(.A1(new_n959), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g830(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g831(.A1(new_n967), .A2(new_n965), .ZN(new_n968));
  INV_X1    g832(.A(KEYINPUT61), .ZN(new_n969));
  INV_X1    g833(.A(new_n943), .ZN(new_n970));
  OAI211_X1 g834(.A(new_n969), .B(new_n970), .C1(new_n957), .C2(KEYINPUT62), .ZN(new_n971));
  OAI21_X1  g835(.A(new_n948), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g836(.A1(new_n966), .A2(new_n972), .ZN(G405));
  INV_X1    g837(.A(new_n952), .ZN(new_n974));
  OAI21_X1  g838(.A(new_n956), .B1(new_n929), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g839(.A1(new_n928), .A2(new_n952), .A3(new_n941), .ZN(new_n976));
  NAND2_X1  g840(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g841(.A(new_n948), .ZN(new_n978));
  XNOR2_X1  g842(.A(new_n977), .B(new_n978), .ZN(G402));
endmodule


