//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n206), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G226gat), .A2(G233gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT77), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G169gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n224), .B(new_n225), .C1(new_n227), .C2(KEYINPUT24), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n216), .A3(new_n218), .A4(KEYINPUT66), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n221), .A2(new_n228), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT24), .B1(new_n226), .B2(KEYINPUT67), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(KEYINPUT67), .B2(new_n226), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n224), .A3(new_n225), .ZN(new_n239));
  NOR2_X1   g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n236), .B1(new_n240), .B2(KEYINPUT23), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n235), .A2(new_n236), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n229), .B1(new_n232), .B2(KEYINPUT26), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT69), .A3(KEYINPUT26), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT27), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G183gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n252), .A3(new_n223), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n226), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n212), .B1(new_n243), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n236), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n242), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OR3_X1    g060(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT29), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n211), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n210), .B(new_n258), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT79), .ZN(new_n267));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n212), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n243), .B2(new_n257), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n261), .A2(new_n262), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n270), .A2(new_n272), .B1(new_n273), .B2(new_n264), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n265), .B(new_n269), .C1(new_n274), .C2(new_n210), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n270), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n264), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n210), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n282), .A2(KEYINPUT30), .A3(new_n265), .A4(new_n269), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n269), .B(KEYINPUT80), .ZN(new_n284));
  INV_X1    g083(.A(new_n265), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n210), .B1(new_n278), .B2(new_n279), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n277), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n290));
  XOR2_X1   g089(.A(G127gat), .B(G134gat), .Z(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(KEYINPUT1), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G113gat), .B(G120gat), .Z(new_n294));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302));
  NOR2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT82), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G148gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n308), .A3(G141gat), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(KEYINPUT83), .A3(new_n311), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n304), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n305), .A2(G141gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT2), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n318), .A2(new_n301), .A3(new_n303), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n298), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n304), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n309), .A2(KEYINPUT83), .A3(new_n311), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT83), .B1(new_n309), .B2(new_n311), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n319), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n293), .A2(new_n297), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n290), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n316), .B2(new_n319), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n324), .A2(new_n333), .A3(new_n325), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n334), .A3(new_n298), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT4), .A4(new_n325), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n331), .B1(new_n339), .B2(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n342), .A2(new_n329), .A3(new_n335), .A4(new_n290), .ZN(new_n343));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT0), .ZN(new_n345));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT85), .B(KEYINPUT6), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n348), .A2(KEYINPUT86), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT86), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n340), .B2(new_n343), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n349), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n289), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n316), .A2(new_n319), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n206), .A2(new_n207), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n206), .A2(new_n207), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n271), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n359), .B1(new_n333), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n210), .B1(new_n334), .B2(new_n271), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n358), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n210), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n368), .B2(new_n359), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G22gat), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n365), .B(new_n372), .C1(new_n364), .C2(new_n369), .ZN(new_n373));
  XOR2_X1   g172(.A(G78gat), .B(G106gat), .Z(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT31), .B(G50gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n371), .A2(KEYINPUT87), .A3(new_n373), .A4(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n380), .A2(new_n376), .B1(new_n371), .B2(new_n373), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n261), .A2(new_n262), .A3(new_n326), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n298), .B1(new_n243), .B2(new_n257), .ZN(new_n384));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT64), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT34), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(new_n387), .B2(KEYINPUT73), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n390), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n383), .A2(new_n384), .A3(new_n387), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n387), .B1(new_n383), .B2(new_n384), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n396));
  XOR2_X1   g195(.A(G15gat), .B(G43gat), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT72), .ZN(new_n398));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n395), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n394), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n326), .B1(new_n261), .B2(new_n262), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n243), .A2(new_n257), .A3(new_n298), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n386), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT70), .A3(new_n401), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT70), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n395), .B2(KEYINPUT33), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n412), .A3(KEYINPUT32), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT71), .B1(new_n395), .B2(new_n396), .ZN(new_n414));
  INV_X1    g213(.A(new_n400), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n404), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n403), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n411), .B2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n394), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n382), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT35), .B1(new_n357), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n400), .B1(new_n424), .B2(KEYINPUT71), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n413), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n404), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n420), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n380), .A2(new_n376), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n371), .A2(new_n373), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n377), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n288), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n277), .A2(new_n283), .A3(KEYINPUT88), .A4(new_n287), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n348), .A2(new_n349), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n355), .B1(new_n441), .B2(new_n352), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n431), .A2(new_n436), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n357), .A2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n427), .B2(new_n404), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n420), .A2(new_n447), .A3(KEYINPUT74), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT74), .B1(new_n420), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(KEYINPUT75), .A2(new_n417), .B1(new_n419), .B2(new_n394), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT36), .B1(new_n451), .B2(new_n429), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n445), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n282), .A2(new_n454), .A3(new_n265), .ZN(new_n455));
  INV_X1    g254(.A(new_n269), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n282), .B2(new_n265), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n281), .B(new_n258), .C1(new_n263), .C2(new_n264), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT37), .C1(new_n274), .C2(new_n281), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n455), .A2(new_n460), .A3(new_n284), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n275), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n382), .B1(new_n464), .B2(new_n442), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT90), .B(KEYINPUT39), .Z(new_n467));
  AND3_X1   g266(.A1(new_n339), .A2(KEYINPUT89), .A3(new_n330), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT89), .B1(new_n339), .B2(new_n330), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n332), .A2(new_n334), .A3(new_n298), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n330), .B1(new_n471), .B2(new_n341), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n339), .A2(KEYINPUT89), .A3(new_n330), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n320), .A2(new_n329), .A3(new_n327), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n476), .A2(KEYINPUT39), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n470), .A2(new_n478), .A3(new_n347), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n352), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n470), .A2(new_n478), .A3(KEYINPUT40), .A4(new_n347), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n466), .B1(new_n484), .B2(new_n440), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n438), .A2(new_n439), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n483), .A2(new_n482), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(KEYINPUT91), .A3(new_n481), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n465), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n444), .B1(new_n453), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT92), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n444), .B(new_n492), .C1(new_n453), .C2(new_n489), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G50gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G43gat), .ZN(new_n496));
  INV_X1    g295(.A(G43gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT94), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT15), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT95), .B1(new_n497), .B2(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n498), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n496), .A2(KEYINPUT95), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n508), .A2(KEYINPUT96), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT14), .B(G29gat), .ZN(new_n510));
  INV_X1    g309(.A(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n503), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n503), .B1(new_n508), .B2(KEYINPUT96), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT97), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT97), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G1gat), .B2(new_n525), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G8gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n517), .B2(new_n519), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n521), .A2(new_n523), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT98), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G197gat), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT11), .B(G169gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n529), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n534), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n536), .B(KEYINPUT13), .Z(new_n550));
  AOI22_X1  g349(.A1(new_n537), .A2(new_n538), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n530), .A2(new_n535), .A3(KEYINPUT18), .A4(new_n536), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n551), .B(new_n552), .C1(new_n539), .C2(new_n545), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n494), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n353), .A2(new_n356), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT7), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  INV_X1    g360(.A(G85gat), .ZN(new_n562));
  INV_X1    g361(.A(G92gat), .ZN(new_n563));
  AOI22_X1  g362(.A1(KEYINPUT8), .A2(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n524), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n532), .A2(new_n567), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n534), .B2(KEYINPUT17), .ZN(new_n570));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT104), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G190gat), .B(G218gat), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n575), .A2(new_n576), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n575), .A2(new_n576), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n585), .B2(new_n577), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G64gat), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n591), .A2(G57gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(G57gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n590), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n600));
  NOR2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(new_n588), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n600), .B(new_n603), .C1(new_n602), .C2(new_n588), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT101), .B(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G127gat), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n605), .A2(KEYINPUT102), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n599), .B2(new_n604), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT21), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n623), .A2(KEYINPUT103), .A3(new_n529), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT103), .B1(new_n623), .B2(new_n529), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n299), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n624), .B2(new_n625), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n616), .A2(new_n617), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n617), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n615), .A4(new_n629), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G230gat), .ZN(new_n637));
  INV_X1    g436(.A(G233gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n565), .B(new_n566), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n605), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n567), .A2(new_n599), .A3(new_n604), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT105), .B(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(KEYINPUT10), .B(new_n567), .C1(new_n618), .C2(new_n620), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n639), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n641), .B2(new_n642), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G120gat), .B(G148gat), .Z(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n587), .A2(new_n636), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n557), .A2(new_n558), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g459(.A1(new_n557), .A2(new_n486), .A3(new_n658), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n661), .A2(G8gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT16), .B(G8gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(KEYINPUT42), .B2(new_n664), .ZN(G1325gat));
  NAND2_X1  g465(.A1(new_n557), .A2(new_n658), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT74), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n417), .A2(KEYINPUT36), .ZN(new_n669));
  INV_X1    g468(.A(new_n394), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n427), .B2(new_n418), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n420), .A2(new_n447), .A3(KEYINPUT74), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n430), .A2(new_n446), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n674), .B2(new_n676), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n667), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n430), .A2(G15gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n667), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n382), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(new_n556), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n655), .B(KEYINPUT107), .Z(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n636), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n465), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n483), .A2(new_n482), .ZN(new_n691));
  INV_X1    g490(.A(new_n347), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n474), .A2(new_n475), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n467), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT40), .B1(new_n694), .B2(new_n478), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT91), .B1(new_n696), .B2(new_n486), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n484), .A2(new_n466), .A3(new_n440), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n690), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT106), .B1(new_n450), .B2(new_n452), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n674), .A2(new_n676), .A3(new_n675), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n445), .A4(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n485), .A2(new_n488), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(new_n690), .B1(new_n435), .B2(new_n357), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n679), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n444), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n587), .A2(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n584), .A2(new_n586), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n491), .A2(new_n493), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n689), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n558), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n587), .A2(new_n636), .A3(new_n655), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n494), .A2(new_n556), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n558), .A2(new_n513), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n720), .A2(new_n718), .A3(new_n721), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n717), .A2(new_n722), .A3(new_n723), .ZN(G1328gat));
  OAI21_X1  g523(.A(G36gat), .B1(new_n715), .B2(new_n440), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n486), .A2(new_n511), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT46), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n720), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n431), .A2(new_n497), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n720), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n679), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n734));
  INV_X1    g533(.A(new_n709), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n702), .A2(new_n703), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n679), .A2(new_n706), .A3(KEYINPUT108), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(new_n444), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n733), .B(new_n688), .C1(new_n734), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n732), .B1(new_n740), .B2(G43gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n730), .B1(new_n741), .B2(KEYINPUT109), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n497), .B1(new_n714), .B2(new_n733), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n743), .B(KEYINPUT47), .C1(new_n744), .C2(new_n732), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(G1330gat));
  AOI21_X1  g545(.A(new_n495), .B1(new_n714), .B2(new_n435), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n720), .A2(G50gat), .A3(new_n382), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1331gat));
  AOI22_X1  g551(.A1(new_n736), .A2(new_n737), .B1(new_n422), .B2(new_n443), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n686), .A2(new_n636), .A3(new_n587), .A4(new_n687), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n558), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g556(.A1(new_n753), .A2(new_n440), .A3(new_n754), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  NAND2_X1  g561(.A1(new_n755), .A2(new_n733), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n430), .A2(G71gat), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n763), .A2(G71gat), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n755), .A2(new_n435), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  INV_X1    g567(.A(new_n636), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n686), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n656), .B(new_n770), .C1(new_n710), .C2(new_n713), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n558), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n770), .A2(new_n587), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n753), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n774), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n558), .A2(new_n562), .A3(new_n655), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n772), .A2(new_n562), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  INV_X1    g580(.A(new_n687), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(G92gat), .A3(new_n440), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n778), .A2(new_n783), .B1(KEYINPUT110), .B2(KEYINPUT52), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n770), .A2(new_n656), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n486), .B(new_n785), .C1(new_n734), .C2(new_n739), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  OR2_X1    g586(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n784), .B2(new_n787), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(G1337gat));
  NAND2_X1  g590(.A1(new_n771), .A2(new_n733), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G99gat), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n430), .A2(G99gat), .A3(new_n656), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n779), .B2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n782), .A2(G106gat), .A3(new_n382), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n778), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n435), .B(new_n785), .C1(new_n734), .C2(new_n739), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n657), .A2(new_n556), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n644), .A2(new_n645), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n647), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n644), .A2(new_n645), .A3(new_n639), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n652), .B1(new_n646), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n807), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT112), .A4(KEYINPUT55), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(new_n654), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n554), .B2(new_n555), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n551), .A2(new_n545), .A3(new_n552), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n549), .A2(new_n550), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n536), .B1(new_n530), .B2(new_n535), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n543), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n821), .A2(new_n655), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n587), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n819), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n711), .A2(new_n827), .A3(new_n824), .A4(new_n821), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n806), .B1(new_n829), .B2(new_n769), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n558), .A2(new_n440), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n421), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n556), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n636), .B1(new_n826), .B2(new_n828), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n382), .B1(new_n837), .B2(new_n806), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n831), .A2(new_n430), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n556), .A2(G113gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n836), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  AOI21_X1  g643(.A(G120gat), .B1(new_n835), .B2(new_n655), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n687), .A2(G120gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n842), .B2(new_n846), .ZN(G1341gat));
  NOR3_X1   g646(.A1(new_n841), .A2(new_n610), .A3(new_n769), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n834), .A2(KEYINPUT113), .A3(new_n769), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(G127gat), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT113), .B1(new_n834), .B2(new_n769), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(G1342gat));
  NOR3_X1   g651(.A1(new_n834), .A2(G134gat), .A3(new_n587), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n841), .B2(new_n587), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n814), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT114), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n815), .A3(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n654), .A2(new_n864), .A3(new_n816), .A4(new_n818), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n825), .B1(new_n865), .B2(new_n556), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n828), .B1(new_n866), .B2(new_n711), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n806), .B1(new_n867), .B2(new_n769), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n382), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n860), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n864), .A2(new_n654), .A3(new_n816), .A4(new_n818), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n555), .B2(new_n554), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n587), .B1(new_n874), .B2(new_n825), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n636), .B1(new_n875), .B2(new_n828), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT115), .B(new_n870), .C1(new_n876), .C2(new_n806), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n869), .B1(new_n830), .B2(new_n382), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n872), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n733), .A2(new_n831), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n556), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G141gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n733), .A2(new_n382), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n832), .A2(new_n310), .A3(new_n556), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT117), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT58), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(KEYINPUT117), .B2(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n881), .B2(G141gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n859), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n892), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n886), .B1(G141gat), .B2(new_n881), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n894), .B(KEYINPUT118), .C1(new_n895), .C2(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1344gat));
  OAI21_X1  g696(.A(new_n869), .B1(new_n868), .B2(new_n382), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n870), .B1(new_n837), .B2(new_n806), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n655), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT59), .B(G148gat), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n832), .A2(new_n883), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT59), .B1(new_n904), .B2(new_n656), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n306), .A3(new_n308), .ZN(new_n906));
  INV_X1    g705(.A(new_n879), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n902), .A2(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n903), .B(new_n906), .C1(new_n907), .C2(new_n908), .ZN(G1345gat));
  NOR3_X1   g708(.A1(new_n904), .A2(KEYINPUT119), .A3(new_n769), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(G155gat), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT119), .B1(new_n904), .B2(new_n769), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n879), .A2(new_n880), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n769), .A2(new_n299), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n911), .A2(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1346gat));
  NAND4_X1  g714(.A1(new_n832), .A2(new_n300), .A3(new_n711), .A4(new_n883), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT120), .Z(new_n917));
  NAND3_X1  g716(.A1(new_n879), .A2(new_n711), .A3(new_n880), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G162gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n558), .A2(new_n440), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n830), .A2(new_n421), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(new_n216), .A3(new_n218), .A4(new_n556), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT122), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n839), .A2(new_n431), .A3(new_n925), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n686), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1348gat));
  OAI21_X1  g731(.A(G176gat), .B1(new_n930), .B2(new_n782), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n231), .A3(new_n655), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT123), .ZN(G1349gat));
  OAI21_X1  g735(.A(G183gat), .B1(new_n930), .B2(new_n769), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n927), .A2(new_n250), .A3(new_n252), .A4(new_n636), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n930), .B2(new_n587), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n223), .A3(new_n711), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n945), .B(new_n946), .C1(KEYINPUT61), .C2(new_n944), .ZN(G1351gat));
  NAND2_X1  g746(.A1(new_n679), .A2(new_n925), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n901), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n686), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n830), .A2(new_n948), .A3(new_n382), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n686), .A2(G197gat), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  OAI21_X1  g759(.A(G204gat), .B1(new_n950), .B2(new_n782), .ZN(new_n961));
  INV_X1    g760(.A(G204gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n952), .A2(new_n962), .A3(new_n655), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT62), .Z(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(G1353gat));
  NAND4_X1  g764(.A1(new_n953), .A2(new_n203), .A3(new_n636), .A4(new_n954), .ZN(new_n966));
  INV_X1    g765(.A(new_n948), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n900), .A2(new_n636), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g772(.A(KEYINPUT127), .B(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1354gat));
  OAI21_X1  g774(.A(G218gat), .B1(new_n950), .B2(new_n587), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n955), .A2(new_n204), .A3(new_n711), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1355gat));
endmodule


