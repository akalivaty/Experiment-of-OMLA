//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT68), .B(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n191), .A2(new_n192), .A3(G143), .A4(G214), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT18), .A2(G131), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n204), .B(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n197), .B2(new_n198), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n199), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n195), .A2(new_n209), .A3(new_n196), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n195), .B2(new_n196), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT72), .A3(new_n205), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n205), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT72), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n215), .A3(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n212), .A2(new_n213), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  AND4_X1   g036(.A1(KEYINPUT87), .A2(new_n197), .A3(KEYINPUT17), .A4(G131), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT87), .B1(new_n211), .B2(KEYINPUT17), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n197), .A2(G131), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n195), .A2(new_n209), .A3(new_n196), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n213), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n197), .A2(KEYINPUT17), .A3(G131), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT87), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n217), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n211), .A2(KEYINPUT87), .A3(KEYINPUT17), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n208), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n229), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n229), .A3(new_n240), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT88), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n230), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(G475), .B1(new_n245), .B2(G902), .ZN(new_n246));
  XNOR2_X1  g060(.A(G128), .B(G143), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT90), .ZN(new_n250));
  XOR2_X1   g064(.A(G116), .B(G122), .Z(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(G107), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(KEYINPUT13), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n194), .A2(G128), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n253), .B(G134), .C1(KEYINPUT13), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n247), .B(new_n248), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT14), .A3(G122), .ZN(new_n259));
  OAI211_X1 g073(.A(G107), .B(new_n259), .C1(new_n251), .C2(KEYINPUT14), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n260), .C1(G107), .C2(new_n251), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT70), .B(G217), .Z(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT9), .B(G234), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n263), .A2(G953), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n262), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT15), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G478), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(G234), .A2(G237), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n273), .A2(G952), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n192), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(G902), .A3(new_n273), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n277), .B(KEYINPUT91), .Z(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT21), .B(G898), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT92), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n270), .B1(new_n267), .B2(new_n268), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n272), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n204), .B(KEYINPUT19), .Z(new_n286));
  OAI221_X1 g100(.A(new_n220), .B1(new_n286), .B2(G146), .C1(new_n210), .C2(new_n211), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n229), .B1(new_n240), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n241), .B1(new_n226), .B2(new_n229), .ZN(new_n290));
  INV_X1    g104(.A(new_n242), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G475), .A2(G902), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT89), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n285), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n288), .B1(new_n244), .B2(new_n242), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n297), .A2(KEYINPUT20), .A3(new_n294), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n246), .B(new_n284), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT93), .ZN(new_n300));
  INV_X1    g114(.A(new_n285), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n297), .B2(new_n294), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n292), .A2(new_n295), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(KEYINPUT20), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n246), .A4(new_n284), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G221), .B1(new_n264), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT12), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n228), .B2(G107), .ZN(new_n311));
  INV_X1    g125(.A(G107), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT3), .A3(G104), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G101), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT74), .B1(new_n312), .B2(G104), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n228), .A3(G107), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n228), .A2(G107), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n312), .A2(G104), .ZN(new_n321));
  OAI21_X1  g135(.A(G101), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n194), .A2(G146), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n205), .A2(G143), .ZN(new_n326));
  OAI211_X1 g140(.A(G128), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n205), .A2(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n194), .A2(G146), .ZN(new_n329));
  INV_X1    g143(.A(G128), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n329), .C1(KEYINPUT1), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n323), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n327), .A2(new_n331), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n319), .A4(new_n322), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n323), .A2(new_n332), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT64), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G137), .ZN(new_n343));
  AND2_X1   g157(.A1(KEYINPUT11), .A2(G134), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT11), .A2(G134), .ZN(new_n346));
  NOR2_X1   g160(.A1(KEYINPUT11), .A2(G134), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(G137), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n209), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n209), .B1(new_n345), .B2(new_n348), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n309), .B1(new_n339), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n333), .A2(new_n336), .B1(new_n332), .B2(new_n323), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n355), .A2(KEYINPUT12), .A3(new_n352), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n192), .A2(G227), .ZN(new_n358));
  XOR2_X1   g172(.A(G110), .B(G140), .Z(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n319), .A2(new_n364), .A3(new_n322), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n332), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT0), .A4(G128), .ZN(new_n369));
  XNOR2_X1  g183(.A(G143), .B(G146), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G128), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n316), .A2(new_n318), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n315), .B1(new_n373), .B2(new_n314), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n375));
  AOI21_X1  g189(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n311), .A2(new_n313), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n316), .A2(new_n318), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n319), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n368), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT10), .B1(new_n333), .B2(new_n336), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n362), .B1(new_n384), .B2(new_n352), .ZN(new_n385));
  NOR4_X1   g199(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT78), .A4(new_n353), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n357), .B(new_n361), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n362), .A3(new_n352), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n319), .A2(new_n364), .A3(new_n322), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n364), .B1(new_n319), .B2(new_n322), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n391), .A2(new_n367), .B1(new_n380), .B2(new_n376), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n337), .A2(new_n366), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n352), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n353), .B1(new_n382), .B2(new_n383), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(new_n353), .C1(new_n382), .C2(new_n383), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n388), .A2(new_n395), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n387), .B1(new_n400), .B2(new_n361), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n401), .A2(new_n402), .A3(new_n268), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n357), .B1(new_n385), .B2(new_n386), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n360), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n388), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n399), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n361), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(G469), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n402), .A2(new_n268), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n308), .B1(new_n403), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n372), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(new_n202), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n416), .A2(new_n417), .B1(new_n202), .B2(new_n332), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT82), .B1(new_n415), .B2(new_n202), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G224), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(G953), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n420), .B(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n258), .A2(G119), .ZN(new_n424));
  INV_X1    g238(.A(G119), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT66), .B1(new_n425), .B2(G116), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n258), .A3(G119), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(G113), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT5), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT2), .B(G113), .Z(new_n434));
  AOI22_X1  g248(.A1(new_n430), .A2(new_n433), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n363), .A2(new_n365), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n429), .B(new_n434), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n374), .A2(new_n375), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n380), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n440), .A2(KEYINPUT81), .A3(new_n441), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n441), .B1(new_n440), .B2(new_n443), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n436), .A2(new_n439), .A3(new_n442), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n423), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(new_n421), .B2(G953), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n418), .A2(new_n419), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n420), .A2(new_n455), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n442), .B(KEYINPUT8), .Z(new_n461));
  INV_X1    g275(.A(new_n435), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n323), .A2(KEYINPUT83), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n323), .A2(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n435), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n460), .A2(new_n451), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(G902), .B1(new_n459), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G210), .B1(G237), .B2(G902), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT85), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n454), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n454), .B2(new_n469), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n414), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n413), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n307), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n437), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n341), .A2(new_n343), .A3(new_n248), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n209), .B1(G134), .B2(G137), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(KEYINPUT65), .A3(new_n481), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n334), .A2(new_n349), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n415), .B1(new_n350), .B2(new_n351), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n248), .B2(new_n340), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT64), .B(G137), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n248), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n349), .B1(new_n492), .B2(KEYINPUT65), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n331), .A3(new_n327), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n345), .A2(new_n348), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G131), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n372), .B1(new_n497), .B2(new_n349), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT30), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n486), .A2(new_n487), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n489), .B1(new_n502), .B2(new_n437), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n191), .A2(new_n192), .A3(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT27), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G101), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT29), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n488), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n486), .A2(new_n487), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n437), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n486), .A2(new_n487), .A3(new_n479), .A4(KEYINPUT28), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n507), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n268), .B1(new_n508), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n519), .A3(new_n488), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(KEYINPUT69), .A3(new_n437), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(KEYINPUT28), .A3(new_n521), .ZN(new_n522));
  AND4_X1   g336(.A1(KEYINPUT29), .A2(new_n522), .A3(new_n507), .A4(new_n511), .ZN(new_n523));
  OAI21_X1  g337(.A(G472), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT30), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n500), .B1(new_n486), .B2(new_n487), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n437), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n507), .A3(new_n488), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT31), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n503), .A2(new_n530), .A3(new_n507), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n515), .A2(new_n516), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NOR2_X1   g348(.A1(G472), .A2(G902), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n524), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n425), .A2(G128), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n330), .A2(KEYINPUT23), .A3(G119), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n425), .A2(G128), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(KEYINPUT23), .ZN(new_n543));
  XOR2_X1   g357(.A(KEYINPUT24), .B(G110), .Z(new_n544));
  XNOR2_X1  g358(.A(G119), .B(G128), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n543), .A2(G110), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n204), .A2(new_n205), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n220), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n545), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n550), .A3(G110), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n543), .B2(G110), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n548), .B1(new_n237), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n543), .A2(G110), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n551), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(new_n217), .A3(new_n221), .A4(new_n549), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n548), .A3(new_n558), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n268), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n560), .A2(KEYINPUT25), .A3(new_n268), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n263), .B1(G234), .B2(new_n268), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n564), .A2(new_n548), .A3(new_n558), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n558), .B1(new_n564), .B2(new_n548), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n571), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n539), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n571), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n568), .B2(new_n569), .ZN(new_n580));
  INV_X1    g394(.A(new_n577), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n580), .A2(KEYINPUT73), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n538), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n478), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  INV_X1    g401(.A(new_n583), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n533), .A2(new_n268), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(G472), .B1(new_n533), .B2(new_n535), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n413), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n454), .A2(new_n469), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n471), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n473), .ZN(new_n596));
  INV_X1    g410(.A(new_n414), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n475), .B2(KEYINPUT94), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n281), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n246), .B1(new_n296), .B2(new_n298), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n267), .A2(new_n601), .A3(new_n268), .ZN(new_n602));
  NAND2_X1  g416(.A1(G478), .A2(G902), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n267), .B(KEYINPUT33), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n601), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n592), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  INV_X1    g425(.A(new_n246), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n272), .A2(new_n283), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n292), .A2(new_n285), .A3(new_n295), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n302), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT95), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n617), .A3(new_n302), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n612), .B(new_n613), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n599), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n592), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n312), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT96), .B(KEYINPUT35), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  XNOR2_X1  g438(.A(new_n555), .B(KEYINPUT97), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n580), .B1(new_n627), .B2(new_n576), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n591), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n478), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  NAND2_X1  g446(.A1(new_n596), .A2(new_n598), .ZN(new_n633));
  INV_X1    g447(.A(new_n628), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n538), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n413), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n275), .B1(new_n278), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n619), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XOR2_X1   g455(.A(new_n638), .B(KEYINPUT39), .Z(new_n642));
  OAI211_X1 g456(.A(new_n308), .B(new_n642), .C1(new_n403), .C2(new_n412), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT40), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n474), .A2(new_n475), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT38), .ZN(new_n646));
  INV_X1    g460(.A(new_n613), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n600), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n503), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n507), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n520), .A2(new_n521), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n650), .B(new_n268), .C1(new_n507), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G472), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n536), .B2(new_n537), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n414), .A3(new_n628), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n644), .A2(new_n646), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT98), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  AOI21_X1  g472(.A(new_n605), .B1(new_n304), .B2(new_n246), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n639), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n600), .A2(new_n606), .A3(new_n639), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n413), .A2(new_n635), .ZN(new_n664));
  INV_X1    g478(.A(new_n633), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n661), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  INV_X1    g481(.A(new_n387), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n361), .B1(new_n406), .B2(new_n407), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n268), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n401), .A2(new_n402), .A3(new_n268), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n308), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n584), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n608), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT100), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n608), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND3_X1  g495(.A1(new_n619), .A2(new_n620), .A3(new_n674), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NOR2_X1   g497(.A1(new_n633), .A2(new_n673), .ZN(new_n684));
  INV_X1    g498(.A(new_n635), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n307), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n307), .A2(new_n684), .A3(new_n688), .A4(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND4_X1  g505(.A1(new_n600), .A2(new_n596), .A3(new_n647), .A4(new_n598), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n529), .A2(new_n531), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n507), .B1(new_n522), .B2(new_n511), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n535), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n535), .C1(new_n693), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT103), .B(G472), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n589), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n580), .A2(new_n581), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n589), .A2(KEYINPUT104), .A3(new_n700), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n699), .A2(new_n703), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n671), .A2(new_n281), .A3(new_n308), .A4(new_n672), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n692), .A2(new_n706), .A3(new_n707), .A4(KEYINPUT105), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n706), .A2(new_n707), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n600), .A2(new_n596), .A3(new_n647), .A4(new_n598), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  AND4_X1   g528(.A1(new_n634), .A2(new_n699), .A3(new_n703), .A4(new_n705), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n661), .A2(new_n663), .A3(new_n684), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT106), .B(G125), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n474), .A2(new_n597), .A3(new_n475), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n408), .A2(KEYINPUT107), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n400), .A2(new_n722), .A3(new_n361), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n723), .A3(G469), .A4(new_n405), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n672), .A3(new_n411), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n720), .A2(new_n725), .A3(new_n308), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n661), .A2(new_n726), .A3(new_n663), .A4(new_n585), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n661), .A2(new_n663), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n720), .A2(new_n725), .A3(KEYINPUT42), .A4(new_n308), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n538), .A2(new_n730), .A3(new_n704), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n538), .A2(new_n704), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n719), .A2(new_n727), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n209), .ZN(G33));
  AND2_X1   g550(.A1(new_n726), .A2(new_n585), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n612), .B1(new_n616), .B2(new_n618), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(new_n647), .A3(new_n639), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NAND3_X1  g555(.A1(new_n304), .A2(new_n246), .A3(new_n606), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT43), .Z(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n591), .A3(new_n634), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n720), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n405), .A2(new_n408), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n402), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n721), .A2(new_n723), .A3(KEYINPUT45), .A4(new_n405), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n410), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n672), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n308), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n642), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n748), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  OR2_X1    g575(.A1(new_n758), .A2(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n663), .A2(new_n661), .ZN(new_n765));
  INV_X1    g579(.A(new_n720), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n765), .A2(new_n538), .A3(new_n583), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n764), .A2(KEYINPUT109), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  INV_X1    g587(.A(new_n582), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT73), .B1(new_n580), .B2(new_n581), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n590), .A2(new_n774), .A3(new_n775), .A4(new_n281), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n413), .A2(new_n776), .A3(new_n476), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n613), .A2(KEYINPUT112), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n272), .B2(new_n283), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n304), .A2(new_n246), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n778), .B1(new_n607), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n659), .A2(KEYINPUT111), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n777), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n307), .B(new_n477), .C1(new_n585), .C2(new_n629), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n682), .B1(new_n708), .B2(new_n712), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n608), .A2(new_n677), .A3(new_n674), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n677), .B1(new_n608), .B2(new_n674), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n797), .A3(new_n690), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n661), .A2(new_n726), .A3(new_n663), .A4(new_n715), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n782), .A2(new_n638), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n664), .A2(new_n738), .A3(new_n720), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT42), .B1(new_n728), .B2(new_n737), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n733), .A2(new_n731), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n765), .A2(new_n805), .A3(new_n729), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n803), .B(new_n740), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n713), .A2(new_n690), .A3(new_n679), .A4(new_n682), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n740), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n735), .A2(new_n811), .A3(new_n802), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n812), .A3(new_n813), .A4(new_n792), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n636), .B1(new_n728), .B2(new_n739), .ZN(new_n815));
  INV_X1    g629(.A(new_n308), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n634), .A2(new_n816), .A3(new_n638), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n711), .A2(new_n654), .A3(new_n725), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n716), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n640), .A2(new_n716), .A3(new_n666), .A4(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n808), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT113), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT113), .B1(new_n786), .B2(new_n787), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n807), .A2(new_n809), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n823), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n824), .B2(new_n825), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT54), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n823), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n810), .A2(new_n823), .A3(new_n792), .A4(new_n812), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n839), .B2(new_n825), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n832), .B1(new_n830), .B2(new_n823), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(KEYINPUT118), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n743), .A2(new_n275), .ZN(new_n848));
  INV_X1    g662(.A(new_n673), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n646), .A2(new_n597), .A3(new_n849), .ZN(new_n850));
  OR3_X1    g664(.A1(new_n848), .A2(new_n706), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT50), .B1(new_n851), .B2(KEYINPUT119), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(KEYINPUT119), .A3(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n583), .A2(new_n275), .ZN(new_n855));
  OR4_X1    g669(.A1(new_n654), .A2(new_n766), .A3(new_n673), .A4(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(new_n600), .A3(new_n606), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n848), .A2(new_n673), .A3(new_n766), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n715), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n854), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n671), .A2(new_n816), .A3(new_n672), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n762), .A2(KEYINPUT120), .A3(new_n763), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n848), .A2(new_n706), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n766), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n762), .A2(new_n763), .A3(new_n861), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n860), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n854), .A2(new_n859), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n852), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n865), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT51), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n848), .A2(new_n673), .A3(new_n766), .A4(new_n805), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT48), .Z(new_n876));
  OAI211_X1 g690(.A(G952), .B(new_n274), .C1(new_n856), .C2(new_n607), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n863), .B2(new_n684), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n870), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n836), .A2(new_n846), .A3(new_n847), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT121), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n671), .A2(new_n672), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT49), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n704), .A2(new_n308), .A3(new_n414), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n742), .A2(new_n654), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n646), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT110), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(G75));
  NOR2_X1   g709(.A1(new_n192), .A2(G952), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT123), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n842), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(G902), .A3(new_n471), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n423), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n898), .B1(new_n907), .B2(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n844), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n410), .B(KEYINPUT57), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n401), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n899), .A2(G902), .A3(new_n752), .A4(new_n751), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n896), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND4_X1  g730(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n297), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n297), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n896), .ZN(G60));
  NAND3_X1  g734(.A1(new_n836), .A2(new_n846), .A3(new_n847), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n603), .B(KEYINPUT59), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n604), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n911), .A2(new_n604), .A3(new_n922), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n898), .ZN(G63));
  AOI21_X1  g739(.A(KEYINPUT60), .B1(G217), .B2(G902), .ZN(new_n926));
  AND3_X1   g740(.A1(KEYINPUT60), .A2(G217), .A3(G902), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n899), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n573), .B2(new_n574), .ZN(new_n929));
  INV_X1    g743(.A(new_n627), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n929), .B(new_n897), .C1(new_n930), .C2(new_n928), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n279), .B2(new_n421), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n809), .A2(new_n829), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n276), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n903), .B1(G898), .B2(new_n192), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  AOI21_X1  g753(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n643), .A2(new_n766), .A3(new_n584), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n784), .B2(new_n785), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n748), .B2(new_n759), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT125), .Z(new_n946));
  AND2_X1   g760(.A1(new_n815), .A2(new_n716), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n657), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n946), .A2(new_n950), .A3(new_n772), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n192), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n502), .B(new_n286), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n276), .A2(G900), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n772), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n759), .A2(new_n692), .A3(new_n805), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n735), .A2(new_n811), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n760), .A2(new_n959), .A3(new_n960), .A4(new_n947), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n962), .B2(new_n192), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n942), .B1(new_n954), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n955), .B1(new_n951), .B2(new_n192), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n963), .A3(KEYINPUT126), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n941), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n954), .A2(new_n942), .A3(new_n964), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT126), .B1(new_n966), .B2(new_n963), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n970), .A3(new_n940), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  INV_X1    g788(.A(new_n962), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n798), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n649), .A2(new_n507), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n896), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n946), .A2(new_n950), .A3(new_n772), .A4(new_n936), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n650), .B1(new_n979), .B2(new_n974), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI211_X1 g796(.A(KEYINPUT127), .B(new_n650), .C1(new_n979), .C2(new_n974), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n834), .A2(new_n835), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n650), .A2(new_n974), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n985), .A2(new_n977), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n984), .A2(new_n987), .ZN(G57));
endmodule


