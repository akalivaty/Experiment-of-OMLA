//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G116), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n187), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G119), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n189), .B2(new_n192), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n187), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G137), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n202), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT64), .A3(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n215), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n216), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n210), .A2(new_n219), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT30), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n203), .A2(KEYINPUT65), .A3(G134), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n201), .B2(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n203), .A2(G134), .ZN(new_n229));
  OAI211_X1 g043(.A(G131), .B(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT66), .A2(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT66), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n233), .A2(new_n234), .B1(new_n220), .B2(new_n216), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n213), .A2(new_n215), .A3(new_n237), .A4(new_n216), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n209), .B(new_n230), .C1(new_n235), .C2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n224), .A2(new_n225), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n225), .B1(new_n224), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n199), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G237), .A2(G953), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT27), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G101), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n195), .A2(new_n198), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n224), .A2(new_n249), .A3(new_n240), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n243), .A2(KEYINPUT31), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G902), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G472), .ZN(new_n254));
  INV_X1    g068(.A(new_n248), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n223), .A2(new_n219), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n209), .B2(new_n207), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n230), .A2(new_n209), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n233), .A2(new_n234), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n221), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n238), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n199), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n256), .B1(new_n263), .B2(new_n250), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n250), .A2(new_n256), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n255), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n243), .A2(new_n248), .A3(new_n250), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n253), .A2(new_n254), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT68), .B(KEYINPUT32), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n253), .A2(KEYINPUT32), .A3(new_n270), .A4(new_n254), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n263), .A2(new_n250), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT28), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(new_n248), .A3(new_n265), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT30), .B1(new_n258), .B2(new_n262), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n224), .A2(new_n225), .A3(new_n240), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n249), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n250), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n255), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n277), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n252), .B1(new_n277), .B2(new_n278), .ZN(new_n285));
  OAI21_X1  g099(.A(G472), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n273), .A2(new_n274), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT16), .ZN(new_n288));
  INV_X1    g102(.A(G140), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(G125), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(G125), .ZN(new_n293));
  INV_X1    g107(.A(G125), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G140), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT16), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT71), .A4(G125), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n292), .A2(new_n296), .A3(G146), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n295), .ZN(new_n299));
  INV_X1    g113(.A(G110), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT24), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G110), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n301), .B2(new_n303), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n236), .A2(G119), .ZN(new_n308));
  AND2_X1   g122(.A1(KEYINPUT66), .A2(G128), .ZN(new_n309));
  NOR2_X1   g123(.A1(KEYINPUT66), .A2(G128), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n311), .B2(G119), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT23), .B1(new_n236), .B2(G119), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT70), .B1(new_n188), .B2(G128), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n236), .A3(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .A4(new_n232), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G110), .ZN(new_n321));
  OAI221_X1 g135(.A(new_n298), .B1(G146), .B2(new_n299), .C1(new_n313), .C2(new_n321), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n307), .A2(new_n312), .B1(new_n320), .B2(G110), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n292), .A2(new_n296), .A3(new_n297), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n214), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n298), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n323), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n322), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT22), .B(G137), .ZN(new_n331));
  INV_X1    g145(.A(G221), .ZN(new_n332));
  INV_X1    g146(.A(G234), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n332), .A2(new_n333), .A3(G953), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n331), .B(new_n334), .Z(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n322), .B(new_n335), .C1(new_n328), .C2(new_n329), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G217), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(G234), .B2(new_n252), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n252), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT74), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n252), .A3(new_n338), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT25), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n287), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G478), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n191), .A2(G122), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT14), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT94), .ZN(new_n359));
  INV_X1    g173(.A(G122), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G116), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(KEYINPUT14), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n358), .A2(KEYINPUT94), .ZN(new_n364));
  OAI21_X1  g178(.A(G107), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G107), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n357), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n236), .B2(G143), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n212), .A2(KEYINPUT91), .A3(G128), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n231), .A2(G143), .A3(new_n232), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n201), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n201), .B1(new_n371), .B2(new_n372), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n365), .B(new_n367), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT13), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n212), .A2(KEYINPUT91), .A3(G128), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT91), .B1(new_n212), .B2(G128), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT92), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n372), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT13), .B1(new_n369), .B2(new_n370), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n309), .A2(new_n310), .A3(new_n212), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT92), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n369), .A2(KEYINPUT13), .A3(new_n370), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n361), .A2(new_n357), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n367), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n373), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT93), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT93), .ZN(new_n395));
  AOI211_X1 g209(.A(new_n395), .B(new_n392), .C1(new_n387), .C2(G134), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n376), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT9), .B(G234), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n398), .A2(new_n340), .A3(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n376), .B(new_n399), .C1(new_n394), .C2(new_n396), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n356), .B1(new_n403), .B2(new_n252), .ZN(new_n404));
  AOI211_X1 g218(.A(G902), .B(new_n355), .C1(new_n401), .C2(new_n402), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G952), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  INV_X1    g222(.A(G237), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n333), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G953), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n252), .B(new_n412), .C1(G234), .C2(G237), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(G898), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  INV_X1    g231(.A(G104), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(KEYINPUT87), .A2(G143), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT87), .A2(G143), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n409), .A2(new_n412), .A3(G214), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(G214), .A3(new_n244), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n208), .ZN(new_n427));
  XNOR2_X1  g241(.A(G125), .B(G140), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n214), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n420), .A2(new_n421), .B1(new_n244), .B2(G214), .ZN(new_n430));
  NOR2_X1   g244(.A1(KEYINPUT87), .A2(G143), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G131), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n427), .B(new_n429), .C1(new_n426), .C2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT17), .B(G131), .C1(new_n430), .C2(new_n432), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n208), .A3(new_n425), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT17), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n325), .A3(new_n298), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n419), .B(new_n434), .C1(new_n437), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n428), .A2(KEYINPUT19), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n428), .A2(KEYINPUT19), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n214), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n298), .ZN(new_n449));
  INV_X1    g263(.A(new_n298), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n299), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G146), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT88), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n438), .A2(new_n433), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n419), .B1(new_n456), .B2(new_n434), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n443), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n459), .B(KEYINPUT90), .Z(new_n460));
  OAI21_X1  g274(.A(KEYINPUT20), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n456), .A2(new_n434), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n442), .B1(new_n462), .B2(new_n419), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  INV_X1    g278(.A(new_n460), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n437), .A2(new_n441), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n419), .B1(new_n467), .B2(new_n434), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n252), .B1(new_n468), .B2(new_n443), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n461), .A2(new_n466), .B1(G475), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n406), .A2(new_n416), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n412), .A2(G227), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n472), .B(new_n473), .Z(new_n474));
  INV_X1    g288(.A(new_n210), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT3), .B1(new_n418), .B2(G107), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n366), .A3(G104), .ZN(new_n478));
  INV_X1    g292(.A(G101), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n418), .A2(G107), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n418), .A2(G107), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n366), .A2(G104), .ZN(new_n483));
  OAI21_X1  g297(.A(G101), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT77), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n481), .B(new_n484), .C1(new_n238), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n212), .A2(G146), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT1), .ZN(new_n490));
  OAI21_X1  g304(.A(G128), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n485), .A3(new_n238), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT10), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT78), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n481), .A2(new_n484), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n481), .B2(new_n484), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n261), .B2(new_n238), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n494), .A2(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G101), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT76), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT76), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n505), .A3(G101), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n506), .A4(new_n481), .ZN(new_n507));
  INV_X1    g321(.A(new_n503), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n257), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n475), .B1(new_n501), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n492), .A2(new_n485), .A3(new_n238), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n495), .B1(new_n513), .B2(new_n486), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n499), .A2(new_n500), .ZN(new_n515));
  AND4_X1   g329(.A1(new_n475), .A2(new_n511), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n474), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n511), .A2(new_n514), .A3(new_n515), .A4(new_n475), .ZN(new_n518));
  INV_X1    g332(.A(new_n474), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n238), .B(new_n261), .C1(new_n497), .C2(new_n498), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n494), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT12), .B1(new_n521), .B2(new_n210), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(new_n475), .C1(new_n520), .C2(new_n494), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n518), .B(new_n519), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G469), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n252), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT79), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n512), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n518), .A2(KEYINPUT79), .A3(new_n519), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n518), .B1(new_n522), .B2(new_n524), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n474), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(G469), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n527), .A2(new_n252), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n528), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n398), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n332), .B1(new_n541), .B2(new_n252), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT75), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n471), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G214), .B1(G237), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n188), .A2(KEYINPUT67), .A3(G116), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT5), .B(new_n194), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G113), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n551), .A2(new_n553), .B1(new_n197), .B2(new_n187), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n481), .A2(new_n484), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT78), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n481), .A2(new_n484), .A3(new_n496), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n502), .A2(new_n505), .A3(G101), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n505), .B1(new_n502), .B2(G101), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n195), .A2(new_n198), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G122), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n558), .B(new_n565), .C1(new_n562), .C2(new_n563), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT6), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n231), .A2(new_n232), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n570));
  INV_X1    g384(.A(new_n221), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n294), .B(new_n238), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT80), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n261), .A2(KEYINPUT80), .A3(new_n294), .A4(new_n238), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n257), .A2(G125), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT81), .B(G224), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G953), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT82), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n576), .B2(new_n577), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT6), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n564), .A2(new_n584), .A3(new_n566), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n569), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT83), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT83), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n569), .A2(new_n583), .A3(new_n588), .A4(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n555), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n552), .B1(new_n197), .B2(KEYINPUT5), .ZN(new_n592));
  OAI221_X1 g406(.A(new_n591), .B1(new_n496), .B2(KEYINPUT84), .C1(new_n592), .C2(new_n195), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n565), .B(KEYINPUT8), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n556), .A2(KEYINPUT84), .A3(new_n557), .ZN(new_n595));
  INV_X1    g409(.A(new_n554), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT7), .B1(new_n578), .B2(G953), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n576), .A2(new_n577), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n568), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT85), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n576), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT85), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n577), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n598), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n601), .B1(new_n606), .B2(KEYINPUT86), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT86), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n608), .A3(new_n598), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n590), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n590), .A2(new_n610), .A3(new_n612), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n548), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n353), .A2(new_n546), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT95), .B(G101), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G3));
  NAND4_X1  g433(.A1(new_n590), .A2(new_n610), .A3(KEYINPUT96), .A4(new_n612), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n547), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n590), .A2(new_n612), .A3(new_n610), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n612), .B1(new_n590), .B2(new_n610), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n517), .B2(new_n525), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n538), .B1(new_n627), .B2(new_n527), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n543), .B1(new_n628), .B2(new_n537), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n251), .A2(new_n252), .ZN(new_n631));
  OAI21_X1  g445(.A(G472), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n632), .A2(new_n271), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n629), .A2(new_n633), .A3(new_n352), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n354), .A2(G902), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n386), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n380), .A2(new_n372), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(KEYINPUT92), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n201), .B1(new_n639), .B2(new_n382), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n395), .B1(new_n640), .B2(new_n392), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n388), .A2(KEYINPUT93), .A3(new_n393), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n399), .B1(new_n643), .B2(new_n376), .ZN(new_n644));
  INV_X1    g458(.A(new_n402), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT33), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n401), .A2(new_n647), .A3(new_n402), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n636), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT97), .B(G478), .Z(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n403), .B2(new_n252), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n415), .A3(new_n470), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n626), .A2(new_n634), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  OAI211_X1 g471(.A(new_n470), .B(new_n416), .C1(new_n405), .C2(new_n404), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n626), .A2(new_n634), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  AND3_X1   g476(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT25), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT25), .B1(new_n346), .B2(new_n347), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n664), .A3(new_n342), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n336), .A2(KEYINPUT36), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n330), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n330), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n667), .A2(new_n344), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT98), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n348), .A2(new_n349), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n341), .A3(new_n351), .ZN(new_n672));
  INV_X1    g486(.A(new_n669), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n670), .A2(new_n633), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n546), .A2(new_n616), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  AND3_X1   g497(.A1(new_n670), .A2(new_n287), .A3(new_n675), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n470), .B1(new_n405), .B2(new_n404), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n411), .B1(new_n413), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n684), .A2(new_n629), .A3(new_n689), .A4(new_n626), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  NAND2_X1  g505(.A1(new_n614), .A2(new_n615), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n687), .B(new_n696), .Z(new_n697));
  NOR2_X1   g511(.A1(new_n545), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n695), .B1(KEYINPUT40), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n406), .A2(new_n470), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n255), .B1(new_n243), .B2(new_n250), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n252), .B1(new_n275), .B2(new_n248), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n273), .A2(new_n274), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n669), .B1(new_n350), .B2(new_n351), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n547), .A2(new_n701), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n700), .B(new_n707), .C1(KEYINPUT40), .C2(new_n699), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  AND4_X1   g523(.A1(new_n287), .A2(new_n670), .A3(new_n629), .A4(new_n675), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n469), .A2(G475), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n687), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n714), .B(new_n715), .C1(new_n649), .C2(new_n652), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n401), .A2(new_n647), .A3(new_n402), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n647), .B1(new_n401), .B2(new_n402), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n635), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n652), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n714), .A4(new_n715), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n710), .A2(new_n725), .A3(new_n626), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  NOR2_X1   g541(.A1(new_n627), .A2(new_n527), .ZN(new_n728));
  AOI211_X1 g542(.A(G469), .B(G902), .C1(new_n517), .C2(new_n525), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n728), .A2(new_n729), .A3(new_n542), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n287), .A2(new_n352), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n626), .A2(new_n654), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND3_X1  g548(.A1(new_n614), .A2(new_n625), .A3(new_n615), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n620), .A2(new_n547), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n659), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n287), .A2(new_n730), .A3(new_n352), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n191), .ZN(G18));
  NOR4_X1   g554(.A1(new_n714), .A2(new_n404), .A3(new_n405), .A4(new_n415), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n670), .A2(new_n741), .A3(new_n287), .A4(new_n675), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n735), .A2(new_n736), .A3(new_n730), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n188), .ZN(G21));
  NAND3_X1  g559(.A1(new_n735), .A2(new_n736), .A3(new_n701), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n730), .A2(new_n633), .A3(new_n352), .A4(new_n416), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n360), .ZN(G24));
  NAND2_X1  g563(.A1(new_n632), .A2(new_n271), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n706), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n717), .A2(new_n724), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n743), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT103), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n717), .A2(new_n724), .A3(new_n751), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n743), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n622), .A2(new_n623), .A3(new_n548), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n542), .B1(new_n628), .B2(new_n537), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n287), .A3(new_n352), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n717), .A2(new_n724), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n542), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n540), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n692), .A2(new_n548), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n271), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n274), .A3(new_n286), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n352), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n760), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n725), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND3_X1  g590(.A1(new_n768), .A2(new_n689), .A3(new_n353), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n534), .B2(new_n536), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n527), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n534), .A2(KEYINPUT45), .A3(new_n536), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n539), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n729), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n766), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(new_n697), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n761), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n653), .A2(new_n714), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(KEYINPUT106), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n796), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n798), .B(new_n750), .C1(new_n665), .C2(new_n669), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n791), .B(new_n801), .C1(new_n800), .C2(new_n799), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  XNOR2_X1  g617(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n787), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n786), .A2(new_n766), .A3(new_n804), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n764), .A2(new_n792), .A3(new_n287), .A4(new_n352), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND3_X1  g624(.A1(new_n352), .A2(new_n547), .A3(new_n544), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT108), .Z(new_n812));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n728), .A2(new_n729), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT109), .Z(new_n815));
  OAI211_X1 g629(.A(new_n812), .B(new_n793), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT110), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n705), .B1(new_n815), .B2(new_n813), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n695), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT103), .B1(new_n752), .B2(new_n753), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n756), .A2(new_n743), .A3(new_n755), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n735), .A2(new_n736), .A3(new_n705), .A4(new_n701), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n672), .A2(new_n673), .A3(new_n715), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n826), .B2(new_n767), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n762), .A2(new_n706), .A3(KEYINPUT111), .A4(new_n715), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n726), .A2(new_n690), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n820), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n710), .B(new_n626), .C1(new_n725), .C2(new_n689), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n758), .A2(KEYINPUT52), .A3(new_n833), .A4(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n742), .A2(new_n743), .B1(new_n737), .B2(new_n738), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n748), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n685), .B1(new_n653), .B2(new_n470), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n634), .A2(new_n616), .A3(new_n416), .A4(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n732), .A2(new_n839), .A3(new_n617), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n840), .A3(new_n681), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n761), .A2(new_n762), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n670), .A2(new_n287), .A3(new_n629), .A4(new_n675), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n714), .A2(new_n404), .A3(new_n405), .A4(new_n687), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n624), .A2(new_n844), .A3(new_n547), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n756), .A2(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n775), .A2(new_n777), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n835), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT112), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT113), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  INV_X1    g669(.A(new_n831), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(new_n856), .B2(new_n758), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n823), .A2(new_n831), .A3(new_n820), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n852), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n352), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n410), .A3(new_n750), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n798), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n806), .A2(new_n807), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n815), .A2(new_n543), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n792), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n730), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n792), .A2(new_n410), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n798), .A2(new_n751), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT118), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n865), .A2(new_n705), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n470), .A3(new_n653), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n867), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n694), .A2(new_n871), .A3(new_n547), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT114), .ZN(new_n883));
  INV_X1    g697(.A(new_n881), .ZN(new_n884));
  OR3_X1    g698(.A1(new_n884), .A2(new_n867), .A3(KEYINPUT114), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT116), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n883), .A2(new_n885), .A3(new_n890), .A4(new_n887), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT50), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n882), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n879), .B(KEYINPUT51), .C1(new_n892), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n889), .A2(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  INV_X1    g714(.A(new_n879), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n772), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n798), .A2(new_n903), .A3(new_n872), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT48), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(KEYINPUT119), .A3(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n653), .A2(new_n470), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n876), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n408), .C1(new_n743), .C2(new_n867), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n898), .A2(new_n902), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT120), .B1(new_n864), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(G952), .B2(G953), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n864), .A2(new_n913), .A3(KEYINPUT120), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n819), .B1(new_n915), .B2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n412), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n252), .B1(new_n861), .B2(new_n852), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT56), .B1(new_n920), .B2(G210), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n569), .A2(new_n585), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT121), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n583), .Z(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n921), .B2(new_n925), .ZN(G51));
  AND3_X1   g741(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n928), .B2(new_n850), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n863), .A3(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(KEYINPUT122), .B(KEYINPUT54), .C1(new_n928), .C2(new_n850), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n538), .B(KEYINPUT57), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT123), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n936), .A3(new_n932), .A4(new_n933), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n526), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT124), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n920), .A2(new_n781), .A3(new_n780), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n935), .B2(new_n937), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n918), .B1(new_n940), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(new_n458), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n458), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n918), .ZN(G60));
  NAND2_X1  g764(.A1(new_n646), .A2(new_n648), .ZN(new_n951));
  XOR2_X1   g765(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n952));
  NOR2_X1   g766(.A1(new_n354), .A2(new_n252), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n864), .B2(new_n955), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n951), .A2(new_n931), .A3(new_n932), .A4(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n918), .A3(new_n957), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n861), .B2(new_n852), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n667), .A3(new_n668), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n919), .C1(new_n339), .C2(new_n961), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g778(.A(G953), .B1(new_n578), .B2(new_n414), .ZN(new_n965));
  INV_X1    g779(.A(new_n841), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(G953), .ZN(new_n967));
  INV_X1    g781(.A(new_n923), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(G898), .B2(new_n412), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n967), .B(new_n969), .ZN(G69));
  AOI21_X1  g784(.A(new_n412), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n791), .A2(new_n626), .A3(new_n701), .A4(new_n903), .ZN(new_n972));
  AND4_X1   g786(.A1(new_n758), .A2(new_n775), .A3(new_n777), .A4(new_n833), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n802), .A2(new_n972), .A3(new_n809), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n412), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n279), .A2(new_n280), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n452), .A2(new_n444), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT126), .Z(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(G900), .B2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n971), .B1(new_n982), .B2(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n708), .A2(new_n758), .A3(new_n833), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  NAND4_X1  g799(.A1(new_n353), .A2(new_n698), .A3(new_n761), .A4(new_n838), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n802), .A2(new_n985), .A3(new_n809), .A4(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n982), .B1(new_n988), .B2(new_n979), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  OAI221_X1 g804(.A(new_n982), .B1(KEYINPUT127), .B2(new_n971), .C1(new_n988), .C2(new_n979), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G72));
  AND2_X1   g806(.A1(new_n283), .A2(new_n268), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT63), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n918), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n281), .A2(new_n248), .A3(new_n282), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n987), .A2(new_n702), .B1(new_n974), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n998), .B2(new_n841), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n993), .A2(new_n995), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n854), .B2(new_n1000), .ZN(G57));
endmodule


