

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773;

  BUF_X1 U379 ( .A(n728), .Z(n359) );
  XNOR2_X1 U380 ( .A(n614), .B(n613), .ZN(n728) );
  BUF_X1 U381 ( .A(n609), .Z(n358) );
  AND2_X1 U382 ( .A1(n435), .A2(n434), .ZN(n433) );
  AND2_X1 U383 ( .A1(n609), .A2(n628), .ZN(n612) );
  XNOR2_X1 U384 ( .A(n576), .B(n530), .ZN(n609) );
  XNOR2_X1 U385 ( .A(n420), .B(KEYINPUT105), .ZN(n700) );
  AND2_X1 U386 ( .A1(n401), .A2(n697), .ZN(n428) );
  NOR2_X1 U387 ( .A1(G902), .A2(n736), .ZN(n529) );
  XNOR2_X1 U388 ( .A(n395), .B(n524), .ZN(n543) );
  XNOR2_X1 U389 ( .A(n498), .B(KEYINPUT21), .ZN(n710) );
  XNOR2_X1 U390 ( .A(n748), .B(KEYINPUT77), .ZN(n395) );
  XNOR2_X1 U391 ( .A(G143), .B(G104), .ZN(n463) );
  XNOR2_X1 U392 ( .A(n457), .B(G119), .ZN(n486) );
  AND2_X1 U393 ( .A1(n390), .A2(n389), .ZN(n484) );
  XNOR2_X1 U394 ( .A(G128), .B(G110), .ZN(n500) );
  NAND2_X1 U395 ( .A1(G234), .A2(G237), .ZN(n488) );
  NOR2_X2 U396 ( .A1(n692), .A2(n651), .ZN(n694) );
  XOR2_X2 U397 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n372) );
  AND2_X2 U398 ( .A1(n574), .A2(KEYINPUT28), .ZN(n425) );
  XNOR2_X2 U399 ( .A(n402), .B(n453), .ZN(n594) );
  NOR2_X2 U400 ( .A1(n729), .A2(n594), .ZN(n597) );
  NAND2_X2 U401 ( .A1(n601), .A2(n682), .ZN(n559) );
  NAND2_X1 U402 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U403 ( .A1(n428), .A2(n429), .ZN(n437) );
  AND2_X2 U404 ( .A1(n580), .A2(n358), .ZN(n687) );
  XOR2_X1 U405 ( .A(n521), .B(n508), .Z(n755) );
  BUF_X1 U406 ( .A(n361), .Z(n738) );
  XNOR2_X2 U407 ( .A(n569), .B(n568), .ZN(n391) );
  XNOR2_X2 U408 ( .A(n558), .B(KEYINPUT39), .ZN(n601) );
  XNOR2_X2 U409 ( .A(G146), .B(G125), .ZN(n539) );
  XNOR2_X2 U410 ( .A(G116), .B(KEYINPUT3), .ZN(n457) );
  XNOR2_X2 U411 ( .A(n523), .B(G107), .ZN(n748) );
  XNOR2_X2 U412 ( .A(G110), .B(G104), .ZN(n523) );
  XNOR2_X2 U413 ( .A(n382), .B(KEYINPUT108), .ZN(n607) );
  INV_X1 U414 ( .A(G237), .ZN(n389) );
  INV_X2 U415 ( .A(G953), .ZN(n763) );
  NAND2_X1 U416 ( .A1(n615), .A2(n566), .ZN(n569) );
  BUF_X1 U417 ( .A(n615), .Z(n374) );
  XNOR2_X1 U418 ( .A(n458), .B(KEYINPUT0), .ZN(n615) );
  OR2_X2 U419 ( .A1(n576), .A2(n707), .ZN(n631) );
  INV_X1 U420 ( .A(n647), .ZN(n692) );
  NAND2_X1 U421 ( .A1(n391), .A2(n365), .ZN(n382) );
  AND2_X1 U422 ( .A1(n416), .A2(n415), .ZN(n414) );
  AND2_X1 U423 ( .A1(n610), .A2(n571), .ZN(n442) );
  XOR2_X1 U424 ( .A(KEYINPUT66), .B(n644), .Z(n645) );
  XNOR2_X1 U425 ( .A(n527), .B(n522), .ZN(n396) );
  XNOR2_X1 U426 ( .A(n388), .B(KEYINPUT96), .ZN(n387) );
  INV_X1 U427 ( .A(n521), .ZN(n522) );
  XNOR2_X1 U428 ( .A(G119), .B(KEYINPUT95), .ZN(n499) );
  BUF_X1 U429 ( .A(n583), .Z(n360) );
  XNOR2_X1 U430 ( .A(n384), .B(n482), .ZN(n583) );
  XNOR2_X2 U431 ( .A(n440), .B(KEYINPUT45), .ZN(n647) );
  NOR2_X1 U432 ( .A1(n652), .A2(n694), .ZN(n361) );
  BUF_X1 U433 ( .A(n662), .Z(n362) );
  NOR2_X1 U434 ( .A1(n652), .A2(n694), .ZN(n664) );
  XNOR2_X2 U435 ( .A(n456), .B(n552), .ZN(n707) );
  XNOR2_X2 U436 ( .A(n446), .B(n534), .ZN(n749) );
  XNOR2_X2 U437 ( .A(n486), .B(n485), .ZN(n446) );
  XNOR2_X2 U438 ( .A(n631), .B(KEYINPUT111), .ZN(n582) );
  NOR2_X2 U439 ( .A1(n570), .A2(n710), .ZN(n456) );
  XNOR2_X2 U440 ( .A(n515), .B(n514), .ZN(n570) );
  INV_X1 U441 ( .A(G953), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n483), .B(n379), .ZN(n378) );
  XNOR2_X1 U443 ( .A(G146), .B(G131), .ZN(n483) );
  XNOR2_X1 U444 ( .A(n380), .B(G137), .ZN(n379) );
  INV_X1 U445 ( .A(KEYINPUT5), .ZN(n380) );
  XOR2_X1 U446 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n756) );
  XNOR2_X1 U447 ( .A(n756), .B(n451), .ZN(n524) );
  XNOR2_X1 U448 ( .A(KEYINPUT67), .B(G101), .ZN(n451) );
  XNOR2_X1 U449 ( .A(n648), .B(KEYINPUT84), .ZN(n691) );
  NAND2_X1 U450 ( .A1(n419), .A2(n697), .ZN(n418) );
  AND2_X1 U451 ( .A1(n421), .A2(n422), .ZN(n398) );
  NAND2_X1 U452 ( .A1(n739), .A2(n518), .ZN(n384) );
  XNOR2_X1 U453 ( .A(KEYINPUT74), .B(G469), .ZN(n528) );
  BUF_X1 U454 ( .A(n570), .Z(n410) );
  XNOR2_X1 U455 ( .A(G113), .B(KEYINPUT75), .ZN(n485) );
  XNOR2_X1 U456 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n474) );
  XNOR2_X1 U457 ( .A(G116), .B(G107), .ZN(n472) );
  XNOR2_X1 U458 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n466) );
  XNOR2_X1 U460 ( .A(G902), .B(KEYINPUT15), .ZN(n605) );
  XNOR2_X1 U461 ( .A(n579), .B(KEYINPUT104), .ZN(n627) );
  INV_X1 U462 ( .A(G902), .ZN(n518) );
  AND2_X1 U463 ( .A1(n640), .A2(n639), .ZN(n445) );
  NAND2_X1 U464 ( .A1(n484), .A2(G214), .ZN(n388) );
  XNOR2_X1 U465 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n386) );
  XNOR2_X1 U466 ( .A(G113), .B(G122), .ZN(n461) );
  XOR2_X1 U467 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n462) );
  XNOR2_X1 U468 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n538) );
  INV_X1 U469 ( .A(KEYINPUT48), .ZN(n455) );
  XNOR2_X1 U470 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U471 ( .A(KEYINPUT14), .B(KEYINPUT92), .ZN(n489) );
  OR2_X1 U472 ( .A1(n610), .A2(n575), .ZN(n517) );
  INV_X1 U473 ( .A(KEYINPUT36), .ZN(n436) );
  NOR2_X1 U474 ( .A1(G900), .A2(n491), .ZN(n492) );
  XNOR2_X1 U475 ( .A(n452), .B(n450), .ZN(n665) );
  XNOR2_X1 U476 ( .A(n376), .B(n377), .ZN(n452) );
  XNOR2_X1 U477 ( .A(n460), .B(n378), .ZN(n377) );
  XNOR2_X1 U478 ( .A(KEYINPUT24), .B(KEYINPUT76), .ZN(n506) );
  XNOR2_X1 U479 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n467) );
  XOR2_X1 U480 ( .A(G131), .B(G140), .Z(n521) );
  XNOR2_X1 U481 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U482 ( .A(G146), .ZN(n525) );
  NAND2_X1 U483 ( .A1(n413), .A2(n369), .ZN(n412) );
  INV_X1 U484 ( .A(KEYINPUT113), .ZN(n453) );
  XNOR2_X1 U485 ( .A(n684), .B(KEYINPUT103), .ZN(n599) );
  INV_X1 U486 ( .A(n410), .ZN(n551) );
  INV_X1 U487 ( .A(n583), .ZN(n577) );
  XNOR2_X1 U488 ( .A(n469), .B(G475), .ZN(n470) );
  XNOR2_X1 U489 ( .A(n665), .B(KEYINPUT62), .ZN(n666) );
  XNOR2_X1 U490 ( .A(KEYINPUT16), .B(G122), .ZN(n533) );
  XNOR2_X1 U491 ( .A(n385), .B(n481), .ZN(n739) );
  INV_X1 U492 ( .A(KEYINPUT60), .ZN(n403) );
  INV_X1 U493 ( .A(KEYINPUT56), .ZN(n405) );
  AND2_X1 U494 ( .A1(n374), .A2(n368), .ZN(n363) );
  OR2_X1 U495 ( .A1(n578), .A2(n438), .ZN(n364) );
  AND2_X1 U496 ( .A1(n708), .A2(n567), .ZN(n365) );
  AND2_X1 U497 ( .A1(n447), .A2(KEYINPUT47), .ZN(n366) );
  NOR2_X1 U498 ( .A1(n364), .A2(n517), .ZN(n367) );
  AND2_X1 U499 ( .A1(n633), .A2(n632), .ZN(n368) );
  XOR2_X1 U500 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n369) );
  NAND2_X1 U501 ( .A1(n545), .A2(G214), .ZN(n697) );
  INV_X1 U502 ( .A(n697), .ZN(n438) );
  XOR2_X1 U503 ( .A(n654), .B(n653), .Z(n370) );
  XOR2_X1 U504 ( .A(n660), .B(n659), .Z(n371) );
  XOR2_X1 U505 ( .A(n736), .B(n735), .Z(n373) );
  BUF_X1 U506 ( .A(n574), .Z(n718) );
  AND2_X2 U507 ( .A1(n584), .A2(n577), .ZN(n684) );
  XNOR2_X1 U508 ( .A(n394), .B(n757), .ZN(n736) );
  XNOR2_X1 U509 ( .A(n543), .B(n396), .ZN(n394) );
  BUF_X1 U510 ( .A(n585), .Z(n401) );
  OR2_X1 U511 ( .A1(n698), .A2(n419), .ZN(n415) );
  AND2_X1 U512 ( .A1(n608), .A2(n607), .ZN(n375) );
  NAND2_X1 U513 ( .A1(n676), .A2(n627), .ZN(n447) );
  XNOR2_X1 U514 ( .A(n376), .B(n480), .ZN(n385) );
  XNOR2_X1 U515 ( .A(n376), .B(n520), .ZN(n757) );
  XNOR2_X2 U516 ( .A(n536), .B(G134), .ZN(n376) );
  XNOR2_X2 U517 ( .A(n381), .B(G143), .ZN(n536) );
  XNOR2_X2 U518 ( .A(G128), .B(KEYINPUT65), .ZN(n381) );
  NAND2_X1 U519 ( .A1(n608), .A2(n607), .ZN(n625) );
  XNOR2_X1 U520 ( .A(n383), .B(KEYINPUT32), .ZN(n608) );
  NAND2_X1 U521 ( .A1(n391), .A2(n442), .ZN(n383) );
  AND2_X1 U522 ( .A1(n391), .A2(n610), .ZN(n636) );
  NAND2_X1 U523 ( .A1(n392), .A2(n603), .ZN(n648) );
  XNOR2_X1 U524 ( .A(n393), .B(n455), .ZN(n392) );
  NAND2_X1 U525 ( .A1(n444), .A2(n443), .ZN(n393) );
  XNOR2_X1 U526 ( .A(n449), .B(KEYINPUT73), .ZN(n444) );
  XNOR2_X1 U527 ( .A(n397), .B(KEYINPUT78), .ZN(n441) );
  NAND2_X1 U528 ( .A1(n459), .A2(n624), .ZN(n397) );
  XNOR2_X2 U529 ( .A(n622), .B(n621), .ZN(n769) );
  XNOR2_X1 U530 ( .A(n448), .B(n372), .ZN(n443) );
  NAND2_X1 U531 ( .A1(n398), .A2(n423), .ZN(n427) );
  AND2_X1 U532 ( .A1(n399), .A2(n668), .ZN(G54) );
  XNOR2_X1 U533 ( .A(n737), .B(n373), .ZN(n399) );
  XNOR2_X1 U534 ( .A(n400), .B(n670), .ZN(G57) );
  NAND2_X1 U535 ( .A1(n669), .A2(n668), .ZN(n400) );
  NAND2_X1 U536 ( .A1(n598), .A2(n771), .ZN(n448) );
  XNOR2_X2 U537 ( .A(n559), .B(KEYINPUT40), .ZN(n598) );
  NAND2_X1 U538 ( .A1(n427), .A2(n454), .ZN(n402) );
  AND2_X1 U539 ( .A1(n407), .A2(n668), .ZN(G66) );
  XNOR2_X1 U540 ( .A(n561), .B(n560), .ZN(n439) );
  XNOR2_X1 U541 ( .A(n404), .B(n403), .ZN(G60) );
  NAND2_X1 U542 ( .A1(n408), .A2(n668), .ZN(n404) );
  XNOR2_X1 U543 ( .A(n406), .B(n405), .ZN(G51) );
  NAND2_X1 U544 ( .A1(n409), .A2(n668), .ZN(n406) );
  NAND2_X1 U545 ( .A1(n441), .A2(n445), .ZN(n440) );
  XNOR2_X1 U546 ( .A(n663), .B(n362), .ZN(n407) );
  XNOR2_X1 U547 ( .A(n655), .B(n370), .ZN(n408) );
  XNOR2_X1 U548 ( .A(n661), .B(n371), .ZN(n409) );
  NAND2_X1 U549 ( .A1(n411), .A2(n374), .ZN(n617) );
  INV_X1 U550 ( .A(n728), .ZN(n411) );
  NAND2_X1 U551 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U552 ( .A1(n414), .A2(n412), .ZN(n729) );
  OR2_X1 U553 ( .A1(n700), .A2(n438), .ZN(n413) );
  NAND2_X1 U554 ( .A1(n417), .A2(n698), .ZN(n416) );
  NOR2_X1 U555 ( .A1(n700), .A2(n418), .ZN(n417) );
  INV_X1 U556 ( .A(n369), .ZN(n419) );
  AND2_X1 U557 ( .A1(n583), .A2(n584), .ZN(n420) );
  XNOR2_X2 U558 ( .A(n585), .B(n556), .ZN(n698) );
  NAND2_X1 U559 ( .A1(n632), .A2(n426), .ZN(n421) );
  NAND2_X1 U560 ( .A1(n575), .A2(n426), .ZN(n422) );
  NAND2_X1 U561 ( .A1(n425), .A2(n424), .ZN(n423) );
  INV_X1 U562 ( .A(n575), .ZN(n424) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n426) );
  INV_X1 U564 ( .A(n578), .ZN(n429) );
  NAND2_X1 U565 ( .A1(n517), .A2(n436), .ZN(n434) );
  NAND2_X1 U566 ( .A1(n433), .A2(n430), .ZN(n580) );
  NAND2_X1 U567 ( .A1(n432), .A2(n431), .ZN(n430) );
  NOR2_X1 U568 ( .A1(n517), .A2(n436), .ZN(n431) );
  INV_X1 U569 ( .A(n437), .ZN(n432) );
  NOR2_X2 U570 ( .A1(n439), .A2(n565), .ZN(n458) );
  NOR2_X1 U571 ( .A1(n594), .A2(n439), .ZN(n676) );
  NOR2_X2 U572 ( .A1(G902), .A2(n654), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n446), .B(n524), .ZN(n450) );
  NOR2_X1 U574 ( .A1(n447), .A2(KEYINPUT47), .ZN(n591) );
  NAND2_X1 U575 ( .A1(n593), .A2(n592), .ZN(n449) );
  INV_X1 U576 ( .A(n576), .ZN(n454) );
  INV_X1 U577 ( .A(n707), .ZN(n628) );
  XNOR2_X1 U578 ( .A(n625), .B(KEYINPUT85), .ZN(n459) );
  BUF_X1 U579 ( .A(n608), .Z(n572) );
  AND2_X1 U580 ( .A1(n484), .A2(G210), .ZN(n460) );
  INV_X1 U581 ( .A(KEYINPUT80), .ZN(n590) );
  INV_X1 U582 ( .A(KEYINPUT81), .ZN(n604) );
  XNOR2_X1 U583 ( .A(n691), .B(n604), .ZN(n606) );
  NOR2_X1 U584 ( .A1(n554), .A2(n710), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n466), .B(n465), .ZN(n468) );
  BUF_X1 U586 ( .A(n676), .Z(n680) );
  XNOR2_X1 U587 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U588 ( .A(n539), .B(n467), .ZN(n508) );
  XNOR2_X1 U589 ( .A(n468), .B(n755), .ZN(n654) );
  XNOR2_X1 U590 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n469) );
  XNOR2_X2 U591 ( .A(n471), .B(n470), .ZN(n584) );
  XOR2_X1 U592 ( .A(KEYINPUT101), .B(G122), .Z(n473) );
  XNOR2_X1 U593 ( .A(n473), .B(n472), .ZN(n477) );
  XOR2_X1 U594 ( .A(KEYINPUT102), .B(KEYINPUT100), .Z(n475) );
  XNOR2_X1 U595 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U596 ( .A(n477), .B(n476), .Z(n481) );
  XOR2_X1 U597 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n479) );
  NAND2_X1 U598 ( .A1(G234), .A2(n763), .ZN(n478) );
  XNOR2_X1 U599 ( .A(n479), .B(n478), .ZN(n503) );
  NAND2_X1 U600 ( .A1(G217), .A2(n503), .ZN(n480) );
  INV_X1 U601 ( .A(G478), .ZN(n482) );
  OR2_X1 U602 ( .A1(n584), .A2(n577), .ZN(n578) );
  NAND2_X1 U603 ( .A1(n665), .A2(n518), .ZN(n487) );
  XNOR2_X2 U604 ( .A(n487), .B(G472), .ZN(n574) );
  XNOR2_X1 U605 ( .A(n574), .B(KEYINPUT6), .ZN(n610) );
  NAND2_X1 U606 ( .A1(n493), .A2(G902), .ZN(n490) );
  XNOR2_X1 U607 ( .A(n490), .B(KEYINPUT93), .ZN(n562) );
  NAND2_X1 U608 ( .A1(G953), .A2(n562), .ZN(n491) );
  XOR2_X1 U609 ( .A(KEYINPUT109), .B(n492), .Z(n494) );
  NAND2_X1 U610 ( .A1(G952), .A2(n493), .ZN(n727) );
  NOR2_X1 U611 ( .A1(n727), .A2(G953), .ZN(n563) );
  NOR2_X1 U612 ( .A1(n494), .A2(n563), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n605), .A2(G234), .ZN(n495) );
  XNOR2_X1 U614 ( .A(n495), .B(KEYINPUT20), .ZN(n512) );
  INV_X1 U615 ( .A(n512), .ZN(n497) );
  INV_X1 U616 ( .A(G221), .ZN(n496) );
  OR2_X1 U617 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X2 U618 ( .A(G137), .B(KEYINPUT72), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n519), .B(n499), .ZN(n502) );
  XNOR2_X1 U620 ( .A(n500), .B(G140), .ZN(n501) );
  XNOR2_X1 U621 ( .A(n502), .B(n501), .ZN(n505) );
  NAND2_X1 U622 ( .A1(n503), .A2(G221), .ZN(n504) );
  XNOR2_X1 U623 ( .A(n505), .B(n504), .ZN(n511) );
  XOR2_X1 U624 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n507) );
  XNOR2_X1 U625 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U627 ( .A(n511), .B(n510), .ZN(n662) );
  NAND2_X1 U628 ( .A1(n662), .A2(n518), .ZN(n515) );
  NAND2_X1 U629 ( .A1(n512), .A2(G217), .ZN(n513) );
  XNOR2_X1 U630 ( .A(n513), .B(KEYINPUT25), .ZN(n514) );
  NAND2_X1 U631 ( .A1(n570), .A2(n516), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n518), .A2(n389), .ZN(n545) );
  INV_X1 U633 ( .A(n519), .ZN(n520) );
  NAND2_X1 U634 ( .A1(G227), .A2(n763), .ZN(n526) );
  XNOR2_X2 U635 ( .A(n529), .B(n528), .ZN(n576) );
  INV_X1 U636 ( .A(KEYINPUT1), .ZN(n530) );
  INV_X1 U637 ( .A(n358), .ZN(n708) );
  NAND2_X1 U638 ( .A1(n367), .A2(n708), .ZN(n532) );
  XNOR2_X1 U639 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n531) );
  XNOR2_X1 U640 ( .A(n532), .B(n531), .ZN(n550) );
  XNOR2_X1 U641 ( .A(n533), .B(KEYINPUT79), .ZN(n534) );
  NAND2_X1 U642 ( .A1(n763), .A2(G224), .ZN(n535) );
  XNOR2_X1 U643 ( .A(n535), .B(KEYINPUT87), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n536), .B(n537), .ZN(n541) );
  XNOR2_X1 U645 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U646 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U647 ( .A(n749), .B(n542), .ZN(n544) );
  XNOR2_X1 U648 ( .A(n544), .B(n543), .ZN(n660) );
  INV_X1 U649 ( .A(n605), .ZN(n643) );
  OR2_X2 U650 ( .A1(n660), .A2(n643), .ZN(n548) );
  NAND2_X1 U651 ( .A1(n545), .A2(G210), .ZN(n546) );
  XNOR2_X1 U652 ( .A(n546), .B(KEYINPUT91), .ZN(n547) );
  XNOR2_X2 U653 ( .A(n548), .B(n547), .ZN(n585) );
  INV_X1 U654 ( .A(n401), .ZN(n549) );
  NAND2_X1 U655 ( .A1(n550), .A2(n549), .ZN(n602) );
  XNOR2_X1 U656 ( .A(n602), .B(G140), .ZN(G42) );
  INV_X1 U657 ( .A(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U658 ( .A1(n574), .A2(n697), .ZN(n553) );
  XNOR2_X1 U659 ( .A(n553), .B(KEYINPUT30), .ZN(n555) );
  NOR2_X1 U660 ( .A1(n555), .A2(n554), .ZN(n581) );
  INV_X1 U661 ( .A(KEYINPUT38), .ZN(n556) );
  AND2_X1 U662 ( .A1(n581), .A2(n698), .ZN(n557) );
  NAND2_X1 U663 ( .A1(n582), .A2(n557), .ZN(n558) );
  INV_X1 U664 ( .A(n578), .ZN(n682) );
  XNOR2_X1 U665 ( .A(n598), .B(G131), .ZN(G33) );
  NAND2_X1 U666 ( .A1(n585), .A2(n697), .ZN(n561) );
  INV_X1 U667 ( .A(KEYINPUT19), .ZN(n560) );
  NOR2_X1 U668 ( .A1(G898), .A2(n763), .ZN(n751) );
  AND2_X1 U669 ( .A1(n562), .A2(n751), .ZN(n564) );
  NOR2_X1 U670 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U671 ( .A1(n700), .A2(n710), .ZN(n566) );
  NOR2_X1 U672 ( .A1(n718), .A2(n551), .ZN(n567) );
  XNOR2_X1 U673 ( .A(n607), .B(G110), .ZN(G12) );
  XNOR2_X1 U674 ( .A(G119), .B(KEYINPUT127), .ZN(n573) );
  INV_X1 U675 ( .A(KEYINPUT22), .ZN(n568) );
  XNOR2_X1 U676 ( .A(n410), .B(KEYINPUT106), .ZN(n711) );
  AND2_X1 U677 ( .A1(n358), .A2(n711), .ZN(n571) );
  XOR2_X1 U678 ( .A(n573), .B(n572), .Z(G21) );
  INV_X1 U679 ( .A(n574), .ZN(n632) );
  NAND2_X1 U680 ( .A1(n578), .A2(n599), .ZN(n579) );
  NOR2_X1 U681 ( .A1(n366), .A2(n687), .ZN(n589) );
  AND2_X1 U682 ( .A1(n582), .A2(n581), .ZN(n587) );
  NOR2_X1 U683 ( .A1(n584), .A2(n360), .ZN(n618) );
  AND2_X1 U684 ( .A1(n401), .A2(n618), .ZN(n586) );
  NAND2_X1 U685 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U686 ( .A(KEYINPUT112), .B(n588), .ZN(n772) );
  AND2_X1 U687 ( .A1(n589), .A2(n772), .ZN(n593) );
  XNOR2_X1 U688 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U689 ( .A(KEYINPUT42), .B(KEYINPUT116), .ZN(n595) );
  XNOR2_X1 U690 ( .A(n595), .B(KEYINPUT115), .ZN(n596) );
  XNOR2_X1 U691 ( .A(n597), .B(n596), .ZN(n771) );
  INV_X1 U692 ( .A(n599), .ZN(n600) );
  NAND2_X1 U693 ( .A1(n601), .A2(n600), .ZN(n689) );
  AND2_X1 U694 ( .A1(n602), .A2(n689), .ZN(n603) );
  NOR2_X1 U695 ( .A1(n606), .A2(n605), .ZN(n641) );
  INV_X1 U696 ( .A(n610), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U698 ( .A(KEYINPUT33), .ZN(n613) );
  INV_X1 U699 ( .A(KEYINPUT34), .ZN(n616) );
  XNOR2_X1 U700 ( .A(n617), .B(n616), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n622) );
  INV_X1 U702 ( .A(KEYINPUT82), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT35), .ZN(n621) );
  INV_X1 U704 ( .A(KEYINPUT44), .ZN(n623) );
  AND2_X1 U705 ( .A1(n769), .A2(n623), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n375), .A2(n769), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n626), .A2(KEYINPUT44), .ZN(n640) );
  INV_X1 U708 ( .A(n627), .ZN(n702) );
  AND2_X1 U709 ( .A1(n358), .A2(n718), .ZN(n629) );
  AND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n720) );
  NAND2_X1 U711 ( .A1(n374), .A2(n720), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT31), .ZN(n685) );
  INV_X1 U713 ( .A(n631), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n685), .A2(n363), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n702), .A2(n634), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n358), .A2(n711), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U718 ( .A(n637), .B(KEYINPUT107), .ZN(n768) );
  NOR2_X1 U719 ( .A1(n638), .A2(n768), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n641), .A2(n647), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT83), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n643), .A2(KEYINPUT2), .ZN(n644) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n652) );
  BUF_X1 U724 ( .A(n648), .Z(n649) );
  INV_X1 U725 ( .A(n649), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n664), .A2(G475), .ZN(n655) );
  XOR2_X1 U728 ( .A(KEYINPUT88), .B(KEYINPUT59), .Z(n653) );
  INV_X1 U729 ( .A(G952), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n656), .A2(G953), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(KEYINPUT90), .ZN(n668) );
  INV_X1 U732 ( .A(n668), .ZN(n742) );
  NAND2_X1 U733 ( .A1(n664), .A2(G210), .ZN(n661) );
  XOR2_X1 U734 ( .A(KEYINPUT86), .B(KEYINPUT54), .Z(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(KEYINPUT55), .ZN(n659) );
  NAND2_X1 U736 ( .A1(n738), .A2(G217), .ZN(n663) );
  XOR2_X1 U737 ( .A(KEYINPUT63), .B(KEYINPUT89), .Z(n670) );
  NAND2_X1 U738 ( .A1(n361), .A2(G472), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(n669) );
  XOR2_X1 U740 ( .A(G104), .B(KEYINPUT117), .Z(n672) );
  NAND2_X1 U741 ( .A1(n363), .A2(n682), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G6) );
  XOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n674) );
  NAND2_X1 U744 ( .A1(n363), .A2(n684), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U746 ( .A(G107), .B(n675), .ZN(G9) );
  XOR2_X1 U747 ( .A(KEYINPUT29), .B(KEYINPUT118), .Z(n678) );
  NAND2_X1 U748 ( .A1(n680), .A2(n684), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U750 ( .A(G128), .B(n679), .ZN(G30) );
  NAND2_X1 U751 ( .A1(n680), .A2(n682), .ZN(n681) );
  XNOR2_X1 U752 ( .A(n681), .B(G146), .ZN(G48) );
  NAND2_X1 U753 ( .A1(n685), .A2(n682), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n683), .B(G113), .ZN(G15) );
  NAND2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n686), .B(G116), .ZN(G18) );
  XNOR2_X1 U757 ( .A(n687), .B(G125), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n688), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U759 ( .A(n689), .B(G134), .ZN(n690) );
  XNOR2_X1 U760 ( .A(KEYINPUT120), .B(n690), .ZN(G36) );
  BUF_X1 U761 ( .A(n691), .Z(n759) );
  NOR2_X1 U762 ( .A1(n692), .A2(n759), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n693), .A2(KEYINPUT2), .ZN(n695) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(G953), .A2(n696), .ZN(n733) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U770 ( .A(KEYINPUT123), .B(n705), .Z(n706) );
  NOR2_X1 U771 ( .A1(n359), .A2(n706), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U773 ( .A(n709), .B(KEYINPUT50), .ZN(n716) );
  AND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n714) );
  XOR2_X1 U775 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n712) );
  XNOR2_X1 U776 ( .A(KEYINPUT49), .B(n712), .ZN(n713) );
  XNOR2_X1 U777 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U781 ( .A(KEYINPUT51), .B(n721), .Z(n722) );
  NOR2_X1 U782 ( .A1(n729), .A2(n722), .ZN(n723) );
  NOR2_X1 U783 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U784 ( .A(n725), .B(KEYINPUT52), .ZN(n726) );
  NOR2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n731) );
  NOR2_X1 U786 ( .A1(n729), .A2(n359), .ZN(n730) );
  NOR2_X1 U787 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U789 ( .A(KEYINPUT53), .B(n734), .Z(G75) );
  NAND2_X1 U790 ( .A1(n738), .A2(G469), .ZN(n737) );
  XOR2_X1 U791 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n735) );
  NAND2_X1 U792 ( .A1(n738), .A2(G478), .ZN(n741) );
  XOR2_X1 U793 ( .A(KEYINPUT124), .B(n739), .Z(n740) );
  XNOR2_X1 U794 ( .A(n741), .B(n740), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n743), .A2(n742), .ZN(G63) );
  NAND2_X1 U796 ( .A1(n647), .A2(n763), .ZN(n747) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U799 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n754) );
  XOR2_X1 U801 ( .A(G101), .B(n748), .Z(n750) );
  XOR2_X1 U802 ( .A(n750), .B(n749), .Z(n752) );
  NOR2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(G69) );
  XOR2_X1 U805 ( .A(n756), .B(n755), .Z(n758) );
  XNOR2_X1 U806 ( .A(n757), .B(n758), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n759), .B(n761), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n760), .A2(n763), .ZN(n766) );
  XNOR2_X1 U809 ( .A(n761), .B(G227), .ZN(n762) );
  NOR2_X1 U810 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U811 ( .A1(G900), .A2(n764), .ZN(n765) );
  NAND2_X1 U812 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U813 ( .A(KEYINPUT125), .B(n767), .ZN(G72) );
  XOR2_X1 U814 ( .A(G101), .B(n768), .Z(G3) );
  XNOR2_X1 U815 ( .A(n769), .B(G122), .ZN(n770) );
  XNOR2_X1 U816 ( .A(n770), .B(KEYINPUT126), .ZN(G24) );
  XNOR2_X1 U817 ( .A(G137), .B(n771), .ZN(G39) );
  XOR2_X1 U818 ( .A(n772), .B(G143), .Z(n773) );
  XNOR2_X1 U819 ( .A(KEYINPUT119), .B(n773), .ZN(G45) );
endmodule

