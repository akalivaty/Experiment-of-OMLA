//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G57gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G64gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(G64gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT92), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n210), .A2(new_n206), .A3(G64gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G64gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G57gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT9), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n202), .A3(new_n203), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G127gat), .B(G155gat), .Z(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT94), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n222), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G183gat), .B(G211gat), .Z(new_n226));
  XOR2_X1   g025(.A(new_n225), .B(new_n226), .Z(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(G1gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT89), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n229), .B1(new_n233), .B2(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(new_n217), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n225), .B(new_n226), .ZN(new_n245));
  INV_X1    g044(.A(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G134gat), .B(G162gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT97), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT96), .B(KEYINPUT7), .ZN(new_n253));
  INV_X1    g052(.A(G85gat), .ZN(new_n254));
  INV_X1    g053(.A(G92gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n253), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(KEYINPUT8), .A2(new_n258), .B1(new_n254), .B2(new_n255), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G99gat), .B(G106gat), .Z(new_n261));
  OR2_X1    g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n261), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G36gat), .ZN(new_n266));
  AND2_X1   g065(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G29gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n272), .A2(KEYINPUT15), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(KEYINPUT15), .ZN(new_n274));
  XNOR2_X1  g073(.A(G43gat), .B(G50gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n274), .A2(new_n275), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G232gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n265), .A2(new_n278), .B1(KEYINPUT41), .B2(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n278), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT17), .B1(new_n278), .B2(KEYINPUT88), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n264), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n252), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n284), .A3(new_n252), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n251), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n280), .A2(KEYINPUT41), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT95), .ZN(new_n291));
  XNOR2_X1  g090(.A(G190gat), .B(G218gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n287), .A3(new_n251), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n293), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n286), .A2(new_n287), .A3(new_n251), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(new_n288), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n249), .A2(new_n300), .A3(KEYINPUT98), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT98), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n299), .B2(new_n248), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n263), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n260), .A2(new_n261), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n217), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT99), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n264), .A2(KEYINPUT99), .A3(new_n217), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n263), .A2(KEYINPUT100), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT100), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n260), .A2(new_n315), .A3(new_n261), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n314), .A2(new_n262), .A3(new_n218), .A4(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n265), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n306), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(new_n312), .A3(new_n317), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n306), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G120gat), .B(G148gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G176gat), .B(G204gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  OR2_X1    g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n319), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n305), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n321), .A2(new_n306), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n332), .ZN(new_n333));
  OR2_X1    g132(.A1(G127gat), .A2(G134gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT69), .B(G127gat), .Z(new_n336));
  INV_X1    g135(.A(G134gat), .ZN(new_n337));
  OAI221_X1 g136(.A(new_n334), .B1(new_n335), .B2(KEYINPUT1), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n339));
  INV_X1    g138(.A(G113gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G113gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n343), .A3(G120gat), .ZN(new_n344));
  INV_X1    g143(.A(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G113gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n339), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n339), .A3(new_n346), .ZN(new_n349));
  NAND2_X1  g148(.A1(G127gat), .A2(G134gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT72), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n350), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT1), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n348), .A2(new_n349), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT65), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT23), .B1(new_n362), .B2(KEYINPUT64), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n364), .B(new_n365), .C1(G169gat), .C2(G176gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(G183gat), .A3(G190gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G183gat), .B(G190gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n356), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT66), .B(new_n356), .C1(new_n367), .C2(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n361), .A2(new_n363), .A3(KEYINPUT25), .A4(new_n366), .ZN(new_n377));
  INV_X1    g176(.A(G183gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G183gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n368), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n369), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT67), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT67), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n369), .C1(new_n370), .C2(new_n368), .ZN(new_n386));
  AOI211_X1 g185(.A(KEYINPUT68), .B(new_n377), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n386), .ZN(new_n389));
  INV_X1    g188(.A(new_n377), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n376), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT27), .B(G183gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n380), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT28), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT26), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n362), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n361), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n338), .B(new_n355), .C1(new_n392), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n387), .A2(new_n391), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n374), .A2(new_n375), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n349), .A2(new_n354), .A3(new_n351), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n338), .B1(new_n408), .B2(new_n347), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT34), .ZN(new_n417));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT73), .ZN(new_n419));
  XOR2_X1   g218(.A(G71gat), .B(G99gat), .Z(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  NAND2_X1  g220(.A1(new_n389), .A2(new_n390), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT68), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n389), .A2(new_n388), .A3(new_n390), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n374), .A3(new_n375), .A4(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n425), .A2(new_n409), .A3(new_n402), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n409), .B1(new_n425), .B2(new_n402), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n426), .A2(new_n427), .A3(new_n415), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n421), .B1(new_n428), .B2(KEYINPUT33), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT34), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n430), .A3(new_n415), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n417), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n404), .A2(new_n410), .A3(new_n414), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT32), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n421), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n411), .B2(new_n415), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT34), .B(new_n414), .C1(new_n404), .C2(new_n410), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n432), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n435), .B1(new_n432), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n407), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n402), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT78), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G197gat), .B(G204gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT74), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT22), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n458), .A2(KEYINPUT75), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n458), .A2(KEYINPUT75), .B1(G211gat), .B2(G218gat), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n453), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n460), .ZN(new_n464));
  INV_X1    g263(.A(new_n457), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n454), .A2(new_n455), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT76), .A3(new_n452), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n392), .B2(new_n403), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n425), .A2(KEYINPUT77), .A3(new_n402), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT29), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n451), .B(new_n470), .C1(new_n474), .C2(new_n449), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n449), .A3(new_n473), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n448), .A2(new_n477), .A3(new_n446), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n469), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G8gat), .B(G36gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n481), .B(new_n482), .Z(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n475), .A2(new_n479), .A3(new_n483), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(KEYINPUT30), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n475), .A2(new_n488), .A3(new_n479), .A4(new_n483), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT31), .B(G50gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  AND2_X1   g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(G141gat), .A2(G148gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G155gat), .A2(G162gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT2), .ZN(new_n499));
  NAND2_X1  g298(.A1(G141gat), .A2(G148gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT79), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n502), .A3(new_n500), .ZN(new_n503));
  INV_X1    g302(.A(new_n498), .ZN(new_n504));
  NOR2_X1   g303(.A1(G155gat), .A2(G162gat), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n501), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n500), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(new_n496), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n504), .A2(new_n505), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n499), .B(new_n508), .C1(new_n509), .C2(new_n502), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n467), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT81), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n453), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n467), .A2(new_n512), .A3(new_n452), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n477), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n506), .B2(new_n510), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n477), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n469), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n495), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n511), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n469), .A2(KEYINPUT29), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(KEYINPUT3), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n495), .B1(new_n469), .B2(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n493), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(G22gat), .B1(new_n532), .B2(KEYINPUT82), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n516), .A2(new_n477), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n520), .B1(new_n534), .B2(new_n515), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n524), .B1(new_n535), .B2(new_n511), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n536), .A2(new_n495), .B1(new_n529), .B2(new_n530), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n537), .A2(new_n493), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n539));
  INV_X1    g338(.A(G22gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(new_n540), .C1(new_n537), .C2(new_n493), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n533), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n538), .B1(new_n533), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n511), .B(new_n338), .C1(new_n408), .C2(new_n347), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n506), .A2(KEYINPUT3), .A3(new_n510), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n409), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n511), .A4(new_n338), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G225gat), .A2(G233gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n409), .A2(new_n527), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n554), .B2(new_n545), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT5), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n551), .A2(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n521), .B1(new_n527), .B2(KEYINPUT3), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n558), .A2(new_n409), .B1(new_n545), .B2(new_n546), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(KEYINPUT5), .A3(new_n552), .A4(new_n550), .ZN(new_n560));
  XNOR2_X1  g359(.A(G1gat), .B(G29gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT0), .ZN(new_n562));
  XNOR2_X1  g361(.A(G57gat), .B(G85gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT6), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n557), .B2(new_n560), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT84), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n557), .A2(new_n560), .ZN(new_n572));
  INV_X1    g371(.A(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT84), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n566), .A4(new_n565), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n569), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n444), .A2(new_n490), .A3(new_n544), .A4(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n571), .B1(new_n568), .B2(new_n567), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n490), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n444), .A2(new_n544), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT87), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n444), .A2(new_n585), .A3(new_n544), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n580), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n475), .A2(new_n590), .A3(new_n479), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n451), .B(new_n469), .C1(new_n474), .C2(new_n449), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n476), .A2(new_n470), .A3(new_n478), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT37), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n483), .A2(KEYINPUT38), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n596), .A3(new_n486), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n480), .A2(KEYINPUT37), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT85), .A3(new_n484), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n590), .B1(new_n475), .B2(new_n479), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n483), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n602), .A3(new_n591), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n603), .B2(KEYINPUT38), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n551), .A2(new_n553), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n554), .A2(new_n552), .A3(new_n545), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT39), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n607), .B(new_n573), .C1(KEYINPUT39), .C2(new_n605), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT83), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(KEYINPUT40), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n565), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n610), .B2(new_n608), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n487), .A2(new_n489), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n544), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n443), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n432), .A2(new_n441), .A3(new_n435), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT36), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n442), .A2(new_n443), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n581), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n487), .B2(new_n489), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n618), .A2(new_n620), .B1(new_n622), .B2(new_n544), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n589), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G197gat), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT11), .B(G169gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n239), .B1(new_n282), .B2(new_n283), .ZN(new_n632));
  NAND2_X1  g431(.A1(G229gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n238), .A2(new_n278), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT90), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n631), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n632), .A2(KEYINPUT18), .A3(new_n633), .A4(new_n634), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n238), .B(new_n278), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n633), .B(KEYINPUT13), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n626), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n333), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n621), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  INV_X1    g453(.A(new_n490), .ZN(new_n655));
  INV_X1    g454(.A(new_n333), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n649), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(G8gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT16), .B(G8gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT42), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(KEYINPUT42), .B2(new_n661), .ZN(G1325gat));
  INV_X1    g462(.A(new_n444), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n652), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n616), .A2(KEYINPUT36), .A3(new_n617), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n619), .B1(new_n442), .B2(new_n443), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n652), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(G15gat), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT101), .B(new_n666), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674));
  INV_X1    g473(.A(new_n666), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n652), .B2(new_n670), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(G1326gat));
  INV_X1    g477(.A(new_n544), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n652), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n650), .A2(new_n651), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n332), .A2(new_n248), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n300), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n621), .A2(new_n270), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n615), .B2(new_n623), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n582), .A2(new_n679), .B1(new_n667), .B2(new_n668), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n691), .B(new_n692), .C1(new_n604), .C2(new_n614), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n589), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n299), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n300), .A2(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n696), .A2(new_n697), .B1(new_n626), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n647), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n581), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n703), .A3(new_n704), .ZN(G1328gat));
  NOR2_X1   g504(.A1(new_n490), .A2(G36gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n683), .A2(new_n685), .A3(new_n706), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n702), .B2(new_n490), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G36gat), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n702), .A2(new_n710), .A3(new_n490), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n708), .B(new_n709), .C1(new_n712), .C2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(KEYINPUT104), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n444), .B(new_n685), .C1(new_n657), .C2(new_n649), .ZN(new_n717));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(KEYINPUT104), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n699), .A2(G43gat), .A3(new_n670), .A4(new_n701), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n702), .B2(new_n544), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n544), .A2(G50gat), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT105), .Z(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n686), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(KEYINPUT48), .C1(new_n686), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  NAND4_X1  g531(.A1(new_n301), .A2(new_n700), .A3(new_n331), .A4(new_n303), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT106), .Z(new_n734));
  AND3_X1   g533(.A1(new_n444), .A2(new_n585), .A3(new_n544), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n585), .B1(new_n444), .B2(new_n544), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n622), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT35), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n690), .A2(new_n693), .B1(new_n738), .B2(new_n580), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n621), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g541(.A(new_n490), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n670), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n664), .A2(G71gat), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n749), .A2(G71gat), .B1(new_n740), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n679), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g553(.A1(new_n583), .A2(new_n577), .A3(new_n578), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n737), .A2(KEYINPUT35), .B1(new_n490), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n698), .B1(new_n756), .B2(new_n624), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n249), .A2(new_n647), .A3(new_n332), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n300), .B1(new_n694), .B2(new_n589), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n697), .B1(new_n739), .B2(new_n300), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(KEYINPUT109), .A3(new_n757), .A4(new_n758), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n621), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G85gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n249), .A2(new_n647), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n695), .A2(new_n299), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n759), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n332), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n254), .A3(new_n621), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT110), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n766), .A2(new_n776), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1336gat));
  NOR2_X1   g577(.A1(new_n490), .A2(G92gat), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n760), .A2(new_n781), .A3(new_n490), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n760), .B2(new_n490), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n655), .A3(new_n764), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n786), .A2(G92gat), .B1(new_n772), .B2(new_n779), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G1337gat));
  NAND3_X1  g588(.A1(new_n762), .A2(new_n670), .A3(new_n764), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G99gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n772), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n664), .A2(G99gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(G1338gat));
  NOR2_X1   g593(.A1(new_n544), .A2(G106gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n699), .A2(new_n679), .A3(new_n758), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n799), .B2(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n796), .A2(new_n797), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n762), .A2(new_n679), .A3(new_n764), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n804), .A2(G106gat), .B1(new_n772), .B2(new_n795), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n805), .ZN(G1339gat));
  NAND3_X1  g605(.A1(new_n318), .A2(new_n306), .A3(new_n319), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n318), .A2(KEYINPUT113), .A3(new_n306), .A4(new_n319), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n328), .A3(KEYINPUT54), .A4(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n325), .B1(new_n320), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n330), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT114), .A3(new_n330), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n817), .A2(new_n647), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n637), .A2(new_n631), .A3(new_n640), .A4(new_n643), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n641), .A2(new_n642), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n630), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n331), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n299), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n817), .A2(new_n821), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n299), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n818), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n831), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n248), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n304), .A2(new_n700), .A3(new_n332), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n839), .A3(KEYINPUT116), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n655), .A2(new_n581), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n544), .A3(new_n444), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n700), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n735), .A2(new_n736), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n845), .A2(new_n621), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n845), .A2(new_n853), .A3(new_n621), .A4(new_n850), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n490), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n647), .A2(new_n341), .A3(new_n343), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n848), .B1(new_n855), .B2(new_n856), .ZN(G1340gat));
  NOR3_X1   g656(.A1(new_n847), .A2(new_n345), .A3(new_n332), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n655), .B1(new_n851), .B2(KEYINPUT117), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n331), .A3(new_n854), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n345), .ZN(G1341gat));
  NAND2_X1  g660(.A1(new_n249), .A2(new_n336), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n248), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n855), .A2(new_n862), .B1(new_n336), .B2(new_n863), .ZN(G1342gat));
  NOR2_X1   g663(.A1(new_n300), .A2(G134gat), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT56), .B1(new_n855), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n859), .A2(new_n868), .A3(new_n854), .A4(new_n865), .ZN(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n847), .B2(new_n300), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n846), .A2(new_n669), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n842), .A2(new_n679), .A3(new_n843), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n700), .A2(new_n815), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT55), .B1(new_n819), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n877), .B2(new_n819), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n829), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n300), .ZN(new_n882));
  INV_X1    g681(.A(new_n837), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n249), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND4_X1   g683(.A1(new_n700), .A2(new_n301), .A3(new_n332), .A4(new_n303), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n679), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n872), .B1(new_n875), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(G141gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n700), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n669), .A2(new_n679), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n655), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n845), .A2(new_n621), .A3(new_n647), .A4(new_n893), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n889), .A2(new_n891), .B1(new_n894), .B2(new_n890), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n895), .B2(KEYINPUT120), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(new_n891), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n872), .B(new_n899), .C1(new_n875), .C2(new_n888), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n844), .A2(new_n581), .A3(new_n655), .A4(new_n892), .ZN(new_n901));
  AOI21_X1  g700(.A(G141gat), .B1(new_n901), .B2(new_n647), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n897), .B(new_n898), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n896), .A2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(new_n874), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n842), .A2(new_n679), .A3(new_n843), .A4(new_n905), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n876), .A2(new_n879), .B1(new_n331), .B2(new_n828), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n883), .B1(new_n907), .B2(new_n299), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n885), .B1(new_n908), .B2(new_n248), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n887), .B1(new_n909), .B2(new_n544), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(new_n669), .A3(new_n331), .A4(new_n846), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n889), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n332), .A2(KEYINPUT59), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n901), .B2(new_n331), .ZN(new_n917));
  OAI221_X1 g716(.A(new_n913), .B1(new_n914), .B2(new_n915), .C1(G148gat), .C2(new_n917), .ZN(G1345gat));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n249), .A2(G155gat), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT121), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n889), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(G155gat), .B1(new_n901), .B2(new_n249), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n901), .A2(new_n249), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n922), .B(KEYINPUT122), .C1(new_n926), .C2(G155gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n901), .B2(new_n299), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n299), .A2(G162gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n889), .B2(new_n930), .ZN(G1347gat));
  NOR3_X1   g730(.A1(new_n664), .A2(new_n621), .A3(new_n490), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n845), .A2(new_n544), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n700), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n842), .A2(new_n581), .A3(new_n843), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n849), .A2(new_n490), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n700), .A2(G169gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT123), .ZN(G1348gat));
  INV_X1    g740(.A(G176gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n942), .A3(new_n331), .ZN(new_n943));
  OAI21_X1  g742(.A(G176gat), .B1(new_n933), .B2(new_n332), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  OAI21_X1  g744(.A(G183gat), .B1(new_n933), .B2(new_n248), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n935), .A2(new_n393), .A3(new_n249), .A4(new_n936), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n948), .B(new_n950), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n933), .B2(new_n300), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n380), .A3(new_n299), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  NOR2_X1   g754(.A1(new_n490), .A2(new_n621), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n669), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n906), .B2(new_n910), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n700), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n892), .A2(new_n490), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n935), .A2(new_n647), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(G1352gat));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n842), .A2(new_n581), .A3(new_n843), .A4(new_n962), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n332), .A2(G204gat), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR4_X1   g770(.A1(new_n966), .A2(KEYINPUT125), .A3(KEYINPUT62), .A4(new_n968), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT62), .B1(new_n966), .B2(new_n968), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n332), .B(new_n957), .C1(new_n906), .C2(new_n910), .ZN(new_n975));
  INV_X1    g774(.A(G204gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n972), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n935), .A2(new_n970), .A3(new_n962), .A4(new_n967), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n958), .A2(new_n331), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n982), .A2(new_n983), .A3(new_n985), .A4(new_n974), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n978), .A2(new_n986), .ZN(G1353gat));
  INV_X1    g786(.A(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n988), .B1(new_n958), .B2(new_n249), .ZN(new_n989));
  OR2_X1    g788(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n992), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n249), .A2(new_n988), .ZN(new_n994));
  OAI22_X1  g793(.A1(new_n991), .A2(new_n993), .B1(new_n966), .B2(new_n994), .ZN(G1354gat));
  OAI21_X1  g794(.A(G218gat), .B1(new_n959), .B2(new_n300), .ZN(new_n996));
  OR2_X1    g795(.A1(new_n300), .A2(G218gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n966), .B2(new_n997), .ZN(G1355gat));
endmodule


