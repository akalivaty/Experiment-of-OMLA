//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT73), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(KEYINPUT22), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n206), .B(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n212), .B2(KEYINPUT29), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G141gat), .B(G148gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n214), .B(new_n217), .C1(new_n218), .C2(KEYINPUT2), .ZN(new_n219));
  INV_X1    g018(.A(G141gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n214), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  AOI211_X1 g027(.A(new_n202), .B(new_n203), .C1(new_n213), .C2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n219), .A2(new_n204), .A3(new_n227), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n219), .A2(new_n227), .A3(new_n232), .A4(new_n204), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n212), .ZN(new_n235));
  OR3_X1    g034(.A1(new_n234), .A2(KEYINPUT85), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT85), .B1(new_n234), .B2(new_n235), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n234), .A2(new_n235), .ZN(new_n239));
  INV_X1    g038(.A(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(new_n205), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT29), .B1(new_n211), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n241), .B2(new_n211), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n243), .B2(new_n204), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n239), .A2(new_n244), .B1(new_n202), .B2(new_n203), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT86), .ZN(new_n247));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT84), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT31), .B(G50gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  MUX2_X1   g050(.A(new_n247), .B(new_n246), .S(new_n251), .Z(new_n252));
  AND3_X1   g051(.A1(new_n238), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n238), .B2(new_n245), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n231), .A2(new_n233), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  AND2_X1   g060(.A1(G127gat), .A2(G134gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(G127gat), .A2(G134gat), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(G113gat), .ZN(new_n265));
  INV_X1    g064(.A(G113gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G120gat), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT70), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n257), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n260), .A2(new_n261), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n262), .A2(new_n263), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT70), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n270), .A2(KEYINPUT71), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT69), .B(G127gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n275), .B2(G134gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n265), .A2(new_n267), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n261), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n274), .A2(new_n240), .A3(new_n279), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n269), .A2(new_n273), .B1(new_n278), .B2(new_n276), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n240), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n282), .A2(new_n283), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(KEYINPUT5), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT80), .B1(new_n287), .B2(new_n240), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n280), .A2(new_n228), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n283), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n280), .A2(KEYINPUT80), .A3(new_n228), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n293), .A2(KEYINPUT81), .A3(new_n294), .A4(new_n295), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n298), .A2(KEYINPUT82), .A3(KEYINPUT5), .A4(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n289), .B(KEYINPUT79), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n296), .B2(new_n297), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT82), .B1(new_n304), .B2(new_n299), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n290), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n298), .A2(KEYINPUT5), .A3(new_n299), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(new_n300), .A3(new_n301), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(KEYINPUT88), .A3(new_n290), .ZN(new_n313));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT0), .ZN(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n320));
  AND4_X1   g119(.A1(KEYINPUT4), .A2(new_n274), .A3(new_n240), .A4(new_n279), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT4), .B1(new_n287), .B2(new_n240), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n283), .B1(new_n323), .B2(new_n282), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n294), .B1(new_n293), .B2(new_n295), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT39), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n282), .A2(new_n286), .A3(new_n288), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n326), .A3(new_n294), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n317), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n320), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT40), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n332), .B(new_n333), .C1(new_n327), .C2(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(G183gat), .A3(G190gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G183gat), .B(G190gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n339), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n346), .B2(new_n343), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n338), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(G190gat), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT24), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354));
  INV_X1    g153(.A(new_n343), .ZN(new_n355));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT23), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(KEYINPUT23), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n353), .A2(new_n358), .A3(new_n362), .A4(new_n340), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G226gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n203), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n351), .A2(KEYINPUT27), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G183gat), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n368), .A2(new_n370), .A3(new_n349), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n371), .A2(new_n373), .B1(G183gat), .B2(G190gat), .ZN(new_n374));
  OR2_X1    g173(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n375));
  NAND2_X1  g174(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n359), .A2(new_n361), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n382), .A3(new_n356), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT27), .B(G183gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n349), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n372), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n374), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n364), .A2(new_n367), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n366), .A2(KEYINPUT29), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(new_n364), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n212), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n364), .A2(new_n387), .A3(new_n367), .ZN(new_n392));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n385), .B2(new_n372), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n371), .A2(new_n373), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n396), .A2(new_n383), .B1(new_n363), .B2(new_n348), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n235), .B(new_n392), .C1(new_n397), .C2(new_n389), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n391), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT74), .B(new_n212), .C1(new_n388), .C2(new_n390), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT75), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(KEYINPUT77), .A3(KEYINPUT30), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n400), .B2(new_n401), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n402), .B2(new_n407), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n400), .A2(KEYINPUT76), .A3(new_n406), .A4(new_n401), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n409), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n337), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n255), .B1(new_n319), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n306), .A2(new_n318), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT37), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n391), .A2(new_n398), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n407), .A2(KEYINPUT38), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n424), .A2(new_n425), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n408), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(KEYINPUT89), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n400), .A2(KEYINPUT37), .A3(new_n401), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT90), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n406), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n424), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n433), .B2(new_n406), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT91), .B(KEYINPUT38), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n406), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT90), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n424), .A3(new_n435), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT91), .B1(new_n442), .B2(KEYINPUT38), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n422), .B(new_n432), .C1(new_n439), .C2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n317), .B(new_n290), .C1(new_n302), .C2(new_n305), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n420), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n317), .B1(new_n306), .B2(new_n307), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(new_n313), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n419), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G15gat), .B(G43gat), .Z(new_n450));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n397), .A2(new_n280), .ZN(new_n454));
  INV_X1    g253(.A(G227gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n203), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n364), .A2(new_n387), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n287), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n453), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT34), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n458), .ZN(new_n463));
  INV_X1    g262(.A(new_n456), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT34), .B(new_n456), .C1(new_n454), .C2(new_n458), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n461), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(KEYINPUT32), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n467), .B2(new_n470), .ZN(new_n473));
  AND2_X1   g272(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n474));
  NOR2_X1   g273(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n467), .A2(new_n470), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n468), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n474), .B1(new_n479), .B2(new_n471), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n317), .B1(new_n312), .B2(new_n290), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n422), .B1(new_n446), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n417), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n484), .B2(new_n255), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n472), .A2(new_n473), .A3(new_n255), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n417), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  INV_X1    g288(.A(new_n255), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n479), .A2(new_n489), .A3(new_n490), .A4(new_n471), .ZN(new_n491));
  INV_X1    g290(.A(new_n417), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n422), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n448), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n449), .A2(new_n485), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G113gat), .B(G141gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n501), .B(KEYINPUT12), .Z(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT15), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G43gat), .ZN(new_n508));
  INV_X1    g307(.A(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT15), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n504), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n512), .A3(KEYINPUT95), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT95), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n510), .A2(new_n514), .A3(new_n511), .A4(new_n504), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT14), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT93), .B(G36gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n517), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT94), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT94), .B1(new_n523), .B2(new_n517), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n516), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n507), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(G36gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n518), .A2(KEYINPUT93), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n525), .B(G29gat), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(new_n521), .A3(new_n519), .ZN(new_n534));
  INV_X1    g333(.A(new_n527), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n528), .A2(new_n536), .A3(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n246), .A2(G15gat), .ZN(new_n538));
  INV_X1    g337(.A(G15gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G22gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G1gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(KEYINPUT16), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n538), .A3(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G8gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT97), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n545), .A2(KEYINPUT98), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(KEYINPUT98), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n543), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(new_n553), .A3(G8gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n516), .A2(new_n526), .A3(new_n556), .A4(new_n527), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n559), .A3(new_n557), .ZN(new_n560));
  INV_X1    g359(.A(new_n555), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n537), .B2(new_n557), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n503), .B(new_n558), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n558), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n555), .B1(new_n537), .B2(new_n557), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n503), .B(KEYINPUT13), .Z(new_n569));
  AOI22_X1  g368(.A1(new_n565), .A2(KEYINPUT18), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n502), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(KEYINPUT99), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n564), .A2(new_n575), .A3(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n569), .B1(new_n566), .B2(new_n567), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n578), .B(new_n502), .C1(new_n564), .C2(new_n571), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT100), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n564), .A2(new_n575), .A3(new_n571), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n575), .B1(new_n564), .B2(new_n571), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n584));
  INV_X1    g383(.A(new_n579), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n573), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n496), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n483), .ZN(new_n589));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT7), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n591), .B2(new_n592), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n600), .A3(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n560), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(new_n563), .ZN(new_n607));
  AND2_X1   g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n537), .A2(new_n557), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n605), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n590), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n607), .ZN(new_n620));
  INV_X1    g419(.A(new_n611), .ZN(new_n621));
  INV_X1    g420(.A(new_n590), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n614), .A2(new_n615), .A3(new_n619), .A4(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n625), .A3(new_n612), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT106), .A4(new_n622), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n618), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G71gat), .A2(G78gat), .ZN(new_n631));
  OR2_X1    g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT9), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  INV_X1    g434(.A(G64gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(new_n636), .B2(G57gat), .ZN(new_n637));
  INV_X1    g436(.A(G57gat), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT102), .B1(new_n638), .B2(G64gat), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n636), .A3(G57gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(KEYINPUT101), .A3(G64gat), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n637), .A2(new_n639), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n636), .A2(G57gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n638), .A2(G64gat), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT9), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n632), .A2(new_n631), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n634), .A2(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n555), .B1(KEYINPUT21), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT105), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n648), .A2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G127gat), .B(G155gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT20), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT103), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(G183gat), .B(G211gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n654), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n630), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n599), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n648), .A2(new_n602), .A3(new_n665), .A4(new_n603), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n648), .A2(new_n665), .B1(new_n602), .B2(new_n603), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G230gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n203), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n648), .A2(new_n665), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n604), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT10), .B1(new_n676), .B2(new_n666), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n648), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n677), .A2(new_n679), .B1(new_n670), .B2(new_n203), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n669), .A2(KEYINPUT109), .A3(new_n671), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n674), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n684), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n663), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n588), .A2(new_n589), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g490(.A1(new_n588), .A2(new_n689), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n417), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n550), .B2(new_n693), .ZN(new_n696));
  MUX2_X1   g495(.A(new_n695), .B(new_n696), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g496(.A(new_n481), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n472), .A2(new_n473), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n539), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n692), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n692), .A2(new_n490), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NOR2_X1   g504(.A1(new_n662), .A2(new_n688), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n630), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n588), .A2(new_n517), .A3(new_n589), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n496), .B2(new_n630), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n485), .A2(new_n449), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n488), .A2(new_n495), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n629), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n707), .A2(new_n587), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n483), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n710), .A2(KEYINPUT111), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1328gat));
  NAND2_X1  g523(.A1(new_n588), .A2(new_n708), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n725), .A2(new_n417), .A3(new_n531), .A4(new_n532), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n718), .A2(new_n417), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n523), .B2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n716), .A3(new_n481), .A4(new_n717), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G43gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n700), .A2(new_n508), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n725), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n730), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1330gat));
  NAND4_X1  g536(.A1(new_n712), .A2(new_n716), .A3(new_n255), .A4(new_n717), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n509), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n739), .B2(new_n738), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n588), .A2(new_n509), .A3(new_n255), .A4(new_n708), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(KEYINPUT48), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(G50gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n742), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(G1331gat));
  INV_X1    g547(.A(new_n573), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n581), .A2(new_n579), .A3(new_n582), .A4(KEYINPUT100), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n688), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n663), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n715), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n483), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n638), .ZN(G1332gat));
  INV_X1    g556(.A(new_n755), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n417), .B(KEYINPUT114), .Z(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(KEYINPUT115), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(KEYINPUT115), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n764), .B(new_n766), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n755), .B2(new_n698), .ZN(new_n768));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n700), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n755), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g571(.A1(new_n758), .A2(new_n255), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n752), .A2(new_n662), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n715), .A2(new_n629), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT51), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n715), .A2(new_n778), .A3(new_n629), .A4(new_n775), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n688), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n591), .A3(new_n589), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n712), .A2(new_n716), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n775), .A2(new_n688), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n782), .A2(new_n483), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n591), .B2(new_n784), .ZN(G1336gat));
  NOR2_X1   g584(.A1(new_n759), .A2(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n782), .A2(new_n759), .A3(new_n783), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n787), .B(new_n788), .C1(new_n592), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n783), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n712), .A2(new_n716), .A3(new_n492), .A4(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(G92gat), .ZN(new_n794));
  AND4_X1   g593(.A1(new_n688), .A2(new_n777), .A3(new_n779), .A4(new_n786), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n792), .B2(G92gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n790), .B1(new_n797), .B2(new_n788), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n799), .A3(new_n700), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n782), .A2(new_n698), .A3(new_n783), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(G1338gat));
  XOR2_X1   g601(.A(KEYINPUT117), .B(G106gat), .Z(new_n803));
  NAND3_X1  g602(.A1(new_n712), .A2(new_n716), .A3(new_n791), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n490), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n777), .A2(new_n688), .A3(new_n779), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n490), .A2(G106gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n689), .A2(new_n587), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n562), .A2(new_n563), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n566), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n812), .A2(new_n503), .B1(new_n568), .B2(new_n569), .ZN(new_n813));
  INV_X1    g612(.A(new_n501), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n688), .B(new_n815), .C1(new_n750), .C2(new_n751), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n674), .A2(new_n680), .A3(new_n681), .A4(new_n687), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT10), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n667), .B2(new_n668), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n671), .B1(new_n819), .B2(new_n678), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n687), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n678), .A3(new_n671), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n680), .A2(new_n823), .A3(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n822), .B2(new_n824), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n817), .B(new_n825), .C1(new_n826), .C2(KEYINPUT118), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n825), .A2(new_n817), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n816), .B1(new_n835), .B2(new_n587), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n580), .A2(new_n586), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n815), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n630), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n829), .A2(new_n834), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n836), .A2(new_n630), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n810), .B1(new_n841), .B2(new_n662), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n486), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n759), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n483), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n587), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(new_n266), .ZN(G1340gat));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n753), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(new_n259), .ZN(G1341gat));
  INV_X1    g651(.A(new_n662), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(new_n275), .Z(G1342gat));
  INV_X1    g654(.A(G134gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n630), .A2(new_n492), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n845), .A2(new_n856), .A3(new_n589), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT56), .Z(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n848), .B2(new_n630), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n847), .A2(new_n698), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n842), .A2(new_n255), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n490), .A2(new_n864), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT120), .B1(new_n822), .B2(new_n824), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(KEYINPUT55), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n822), .A2(KEYINPUT120), .A3(new_n824), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n752), .A2(new_n831), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n629), .B1(new_n872), .B2(new_n816), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n838), .A2(new_n835), .A3(new_n630), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n853), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n875), .B2(new_n810), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n862), .B1(new_n865), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n220), .B1(new_n878), .B2(new_n752), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n862), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n752), .A2(new_n220), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT58), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n862), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n842), .B2(new_n255), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  OAI21_X1  g686(.A(G141gat), .B1(new_n887), .B2(new_n587), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n888), .B(new_n889), .C1(new_n881), .C2(new_n882), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n884), .A2(new_n890), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n880), .A2(new_n222), .A3(new_n688), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n827), .A2(new_n828), .ZN(new_n894));
  AND4_X1   g693(.A1(new_n837), .A2(new_n629), .A3(new_n815), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n831), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n816), .B1(new_n587), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n630), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n853), .B1(new_n898), .B2(KEYINPUT121), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n873), .A2(new_n900), .A3(new_n895), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n810), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n255), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n843), .A2(new_n867), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n688), .B(new_n885), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n893), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n222), .C1(new_n878), .C2(new_n688), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n892), .B1(new_n906), .B2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(G155gat), .B1(new_n887), .B2(new_n853), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n880), .A2(new_n215), .A3(new_n662), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1346gat));
  AOI21_X1  g710(.A(new_n216), .B1(new_n878), .B2(new_n629), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n698), .A2(new_n216), .A3(new_n589), .A4(new_n857), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n863), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G162gat), .B1(new_n887), .B2(new_n630), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n916), .B(new_n917), .C1(new_n863), .C2(new_n913), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(G1347gat));
  NAND4_X1  g718(.A1(new_n842), .A2(new_n483), .A3(new_n492), .A4(new_n486), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n840), .A2(new_n752), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n629), .B1(new_n922), .B2(new_n816), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n853), .B1(new_n923), .B2(new_n874), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n589), .B1(new_n924), .B2(new_n810), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n492), .A4(new_n486), .ZN(new_n927));
  AND4_X1   g726(.A1(G169gat), .A2(new_n921), .A3(new_n927), .A4(new_n752), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n486), .A3(new_n846), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n752), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n928), .A2(new_n931), .ZN(G1348gat));
  INV_X1    g731(.A(G176gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n933), .A3(new_n688), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n921), .A2(new_n927), .A3(new_n688), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n933), .ZN(G1349gat));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT125), .Z(new_n939));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n927), .A3(new_n662), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G183gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n842), .A2(new_n483), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n662), .A2(new_n384), .ZN(new_n943));
  NOR4_X1   g742(.A1(new_n942), .A2(new_n844), .A3(new_n759), .A4(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n939), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n939), .ZN(new_n947));
  AOI211_X1 g746(.A(new_n947), .B(new_n944), .C1(new_n940), .C2(G183gat), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n349), .A3(new_n629), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n921), .A2(new_n927), .A3(new_n629), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(G190gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n951), .B2(G190gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n698), .A2(new_n255), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(new_n759), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n942), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n925), .A2(KEYINPUT126), .A3(new_n958), .ZN(new_n961));
  XNOR2_X1  g760(.A(KEYINPUT127), .B(G197gat), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n752), .A4(new_n962), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n903), .A2(new_n904), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n589), .A2(new_n481), .A3(new_n417), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n964), .A2(new_n752), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n966), .B2(new_n962), .ZN(G1352gat));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n688), .A3(new_n965), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G204gat), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n753), .A2(G204gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n925), .A2(new_n958), .A3(new_n970), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT62), .Z(new_n972));
  NAND2_X1  g771(.A1(new_n969), .A2(new_n972), .ZN(G1353gat));
  NAND4_X1  g772(.A1(new_n960), .A2(new_n961), .A3(new_n208), .A4(new_n662), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n662), .B(new_n965), .C1(new_n903), .C2(new_n904), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n961), .A3(new_n209), .A4(new_n629), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n964), .A2(new_n629), .A3(new_n965), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n209), .ZN(G1355gat));
endmodule


