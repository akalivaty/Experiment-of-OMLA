//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  AND2_X1   g0007(.A1(KEYINPUT65), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(KEYINPUT65), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NOR3_X1   g0011(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n212), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n219), .B2(new_n220), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n213), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G107), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n218), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n214), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n222), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(KEYINPUT67), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  OAI21_X1  g0053(.A(G274), .B1(new_n253), .B2(new_n211), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n256), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT67), .A4(G274), .ZN(new_n261));
  INV_X1    g0061(.A(new_n260), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n257), .A2(new_n261), .B1(new_n263), .B2(G226), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT68), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G222), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n277), .B1(new_n229), .B2(new_n275), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n265), .B1(new_n280), .B2(new_n262), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n281), .A2(G169), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT69), .B1(new_n214), .B2(new_n271), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n286), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(new_n211), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n210), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n210), .A2(new_n292), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT70), .A2(G58), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT8), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(new_n271), .A3(KEYINPUT72), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(G20), .B2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n289), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n285), .A2(new_n211), .A3(new_n287), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n255), .A2(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G50), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n305), .A2(new_n307), .B1(G50), .B2(new_n304), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n283), .A2(new_n284), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n311), .ZN(new_n312));
  OR3_X1    g0112(.A1(new_n303), .A2(KEYINPUT9), .A3(new_n308), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT9), .B1(new_n303), .B2(new_n308), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n281), .B2(G190), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT74), .B1(new_n281), .B2(new_n311), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n312), .A2(new_n315), .A3(new_n319), .A4(new_n316), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n310), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n266), .A2(new_n267), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G226), .A2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT80), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n272), .A2(new_n273), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT80), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(G226), .A4(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(G1698), .B1(new_n272), .B2(new_n273), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n262), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n257), .A2(new_n261), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n263), .A2(G232), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(G169), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n260), .B1(new_n328), .B2(new_n330), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n334), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n337), .A2(new_n338), .A3(G179), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT81), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT7), .B1(new_n325), .B2(G20), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n210), .A2(new_n322), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n343), .A3(G68), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n301), .A2(G159), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G58), .A2(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n206), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G20), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT78), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G159), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n298), .B2(new_n300), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n297), .B1(new_n206), .B2(new_n346), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT78), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(KEYINPUT16), .B(new_n344), .C1(new_n349), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n345), .A2(new_n348), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n268), .B1(new_n266), .B2(new_n267), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n273), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT7), .A2(G20), .ZN(new_n360));
  OR2_X1    g0160(.A1(KEYINPUT65), .A2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT65), .A2(G20), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n361), .A2(new_n272), .A3(new_n362), .A4(new_n273), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n359), .A2(new_n360), .B1(KEYINPUT7), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n356), .B1(new_n364), .B2(G68), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n355), .B(new_n288), .C1(new_n365), .C2(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n295), .A2(new_n306), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n367), .A2(new_n305), .B1(new_n304), .B2(new_n295), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n332), .A2(new_n282), .A3(new_n335), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT81), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n337), .B2(new_n338), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n340), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT18), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT18), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n340), .A2(new_n370), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n332), .A2(G190), .A3(new_n335), .ZN(new_n380));
  OAI21_X1  g0180(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n366), .A2(new_n369), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n380), .A2(new_n381), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n366), .A4(new_n369), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n377), .A2(new_n379), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n263), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n333), .B1(new_n230), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n390), .B1(new_n231), .B2(new_n275), .C1(new_n278), .C2(new_n225), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(new_n262), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(G169), .ZN(new_n393));
  XOR2_X1   g0193(.A(KEYINPUT8), .B(G58), .Z(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n301), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT15), .B(G87), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n395), .B1(new_n229), .B2(new_n210), .C1(new_n290), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n288), .ZN(new_n398));
  INV_X1    g0198(.A(new_n305), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n229), .B1(new_n255), .B2(G20), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT73), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n304), .B2(G77), .ZN(new_n402));
  INV_X1    g0202(.A(new_n304), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT73), .A3(new_n229), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n399), .A2(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n393), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n392), .A2(new_n282), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n406), .B1(new_n392), .B2(G190), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n311), .B2(new_n392), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n387), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT76), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n291), .A2(G77), .A3(new_n293), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n301), .A2(G50), .B1(G20), .B2(new_n224), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n289), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .ZN(new_n419));
  OR3_X1    g0219(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n306), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n305), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n418), .A2(KEYINPUT11), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n415), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n418), .B2(KEYINPUT11), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(KEYINPUT76), .C1(KEYINPUT11), .C2(new_n418), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n357), .A2(new_n358), .A3(G226), .A4(new_n276), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n357), .A2(new_n358), .A3(G232), .A4(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G97), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n432), .B(new_n433), .C1(new_n271), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n262), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT75), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n263), .A2(G238), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n333), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n333), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n442));
  INV_X1    g0242(.A(G190), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n436), .B(new_n444), .C1(new_n439), .C2(new_n440), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(G200), .B1(new_n442), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n431), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n333), .A2(new_n438), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n333), .A2(new_n437), .A3(new_n438), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n444), .B1(new_n455), .B2(new_n436), .ZN(new_n456));
  INV_X1    g0256(.A(new_n445), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n311), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n446), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT77), .A3(new_n431), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n431), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n442), .A2(new_n445), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT14), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(G169), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n442), .A2(G179), .A3(new_n445), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n463), .B2(G169), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n321), .A2(new_n414), .A3(new_n461), .A4(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n403), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n271), .A2(G97), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n361), .A2(new_n473), .A3(new_n362), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n297), .A2(G116), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT20), .B1(new_n478), .B2(new_n288), .ZN(new_n479));
  AND4_X1   g0279(.A1(KEYINPUT20), .A2(new_n288), .A3(new_n477), .A4(new_n475), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT89), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n471), .B1(new_n255), .B2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n399), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n483), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT89), .B1(new_n305), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT90), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n478), .A2(KEYINPUT20), .A3(new_n288), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n288), .A2(new_n477), .A3(new_n475), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n484), .A2(new_n486), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT90), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n472), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G41), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n255), .B(G45), .C1(new_n498), .C2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G41), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(KEYINPUT88), .A3(G270), .A4(new_n260), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT88), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n260), .B1(new_n499), .B2(new_n501), .ZN(new_n505));
  INV_X1    g0305(.A(G270), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G303), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n357), .B2(new_n358), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n218), .A2(G1698), .ZN(new_n511));
  OAI221_X1 g0311(.A(new_n511), .B1(G257), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n262), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n254), .ZN(new_n515));
  INV_X1    g0315(.A(new_n499), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n500), .B2(G41), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n515), .A2(new_n516), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n508), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G169), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT21), .B1(new_n497), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(G200), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n443), .B2(new_n521), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n497), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n521), .A2(KEYINPUT21), .A3(G169), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n508), .A2(new_n514), .A3(G179), .A4(new_n520), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n488), .A2(new_n496), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n304), .A2(G97), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n305), .B1(new_n255), .B2(G33), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n231), .A2(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n434), .A2(G107), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT82), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT6), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n536), .A2(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT83), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n361), .A2(new_n362), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT83), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n539), .A2(new_n541), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n544), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n301), .A2(G77), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n360), .B1(new_n269), .B2(new_n274), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n363), .A2(KEYINPUT7), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(G107), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n364), .A2(KEYINPUT85), .A3(G107), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n554), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n535), .B1(new_n563), .B2(new_n289), .ZN(new_n564));
  OAI211_X1 g0364(.A(G244), .B(new_n276), .C1(new_n266), .C2(new_n267), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(G33), .B2(G283), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n357), .A2(new_n358), .A3(G250), .A4(G1698), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n566), .A2(new_n230), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n357), .A2(new_n358), .A3(new_n276), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n262), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n260), .B(G257), .C1(new_n499), .C2(new_n501), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n520), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n373), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n574), .B1(new_n571), .B2(new_n262), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n282), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n564), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n576), .A2(new_n311), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n443), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n535), .B(new_n585), .C1(new_n563), .C2(new_n289), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT22), .B1(new_n275), .B2(G87), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n545), .A2(new_n589), .B1(KEYINPUT23), .B2(G107), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n325), .A2(new_n210), .A3(KEYINPUT22), .A4(G87), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n271), .A2(new_n471), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n297), .B1(new_n592), .B2(KEYINPUT23), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT24), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n590), .A2(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT24), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n359), .B2(new_n226), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n596), .A2(new_n597), .A3(new_n599), .A4(new_n591), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n289), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n534), .A2(G107), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n304), .A2(G107), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT25), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n502), .A2(G264), .A3(new_n260), .ZN(new_n607));
  XOR2_X1   g0407(.A(KEYINPUT91), .B(G294), .Z(new_n608));
  NOR2_X1   g0408(.A1(G250), .A2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n217), .B2(G1698), .ZN(new_n610));
  AOI22_X1  g0410(.A1(G33), .A2(new_n608), .B1(new_n610), .B2(new_n325), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n607), .B(new_n520), .C1(new_n611), .C2(new_n260), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n311), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT92), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT92), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n615), .A3(new_n311), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n612), .A2(G190), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n226), .A2(new_n434), .A3(new_n231), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n621), .A2(new_n271), .A3(new_n434), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n622), .B2(new_n545), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n361), .A2(G33), .A3(G97), .A4(new_n362), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n621), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n325), .A2(new_n210), .A3(G68), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(new_n288), .B1(new_n403), .B2(new_n396), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n534), .A2(G87), .ZN(new_n629));
  INV_X1    g0429(.A(G45), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n213), .B1(new_n630), .B2(G1), .ZN(new_n631));
  INV_X1    g0431(.A(G274), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n255), .A2(new_n632), .A3(G45), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n260), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(G238), .A2(G1698), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n230), .B2(G1698), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n592), .B1(new_n636), .B2(new_n325), .ZN(new_n637));
  OAI211_X1 g0437(.A(G190), .B(new_n634), .C1(new_n637), .C2(new_n260), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n637), .B2(new_n260), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G200), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n628), .A2(new_n629), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n627), .A2(new_n288), .ZN(new_n642));
  INV_X1    g0442(.A(new_n396), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n534), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n396), .A2(new_n403), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(G169), .ZN(new_n647));
  OAI211_X1 g0447(.A(G179), .B(new_n634), .C1(new_n637), .C2(new_n260), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n646), .A2(KEYINPUT87), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT87), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n628), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n641), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n612), .A2(new_n373), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n612), .A2(G179), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(new_n601), .C2(new_n605), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n619), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NOR4_X1   g0456(.A1(new_n470), .A2(new_n532), .A3(new_n587), .A4(new_n656), .ZN(G372));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n318), .A2(new_n320), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n384), .A2(new_n386), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n410), .B1(new_n451), .B2(new_n460), .ZN(new_n662));
  INV_X1    g0462(.A(new_n469), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n377), .A2(new_n379), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n658), .B1(new_n667), .B2(new_n310), .ZN(new_n668));
  INV_X1    g0468(.A(new_n310), .ZN(new_n669));
  INV_X1    g0469(.A(new_n410), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n459), .A2(KEYINPUT77), .A3(new_n431), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT77), .B1(new_n459), .B2(new_n431), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n469), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n665), .B1(new_n674), .B2(new_n661), .ZN(new_n675));
  OAI211_X1 g0475(.A(KEYINPUT93), .B(new_n669), .C1(new_n675), .C2(new_n660), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n470), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n528), .A2(new_n529), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n497), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n522), .B1(new_n488), .B2(new_n496), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n680), .B(new_n655), .C1(KEYINPUT21), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n647), .A2(new_n648), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n646), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n628), .A2(new_n640), .A3(new_n629), .A4(new_n638), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n606), .B2(new_n618), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n682), .A2(new_n582), .A3(new_n586), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n551), .A2(new_n553), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT84), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT85), .B1(new_n364), .B2(G107), .ZN(new_n691));
  INV_X1    g0491(.A(new_n360), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n357), .B2(new_n358), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n342), .B1(new_n210), .B2(new_n322), .ZN(new_n694));
  NOR4_X1   g0494(.A1(new_n693), .A2(new_n694), .A3(new_n558), .A4(new_n231), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n690), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n288), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n580), .B1(new_n699), .B2(new_n535), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n652), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT26), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  INV_X1    g0503(.A(new_n686), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n564), .A2(new_n703), .A3(new_n581), .A4(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n688), .A2(new_n702), .A3(new_n684), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n678), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n677), .A2(new_n707), .ZN(G369));
  NAND3_X1  g0508(.A1(new_n210), .A2(new_n255), .A3(G13), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G213), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(KEYINPUT27), .B2(new_n709), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G343), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n497), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT94), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n524), .A3(new_n530), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n532), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n655), .A2(new_n714), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n619), .B1(new_n606), .B2(new_n713), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n655), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(G330), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT95), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n524), .A2(new_n530), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n714), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n721), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n719), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n729), .ZN(G399));
  NOR2_X1   g0530(.A1(new_n216), .A2(G41), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n255), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n620), .A2(G116), .ZN(new_n733));
  INV_X1    g0533(.A(new_n207), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n731), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n576), .A2(new_n612), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n639), .A2(new_n282), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n521), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n611), .A2(new_n260), .ZN(new_n745));
  INV_X1    g0545(.A(new_n607), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n745), .A2(new_n746), .A3(new_n639), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n578), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n744), .B1(new_n748), .B2(new_n529), .ZN(new_n749));
  INV_X1    g0549(.A(new_n529), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n578), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n714), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT31), .ZN(new_n754));
  INV_X1    g0554(.A(new_n535), .ZN(new_n755));
  AOI221_X4 g0555(.A(new_n755), .B1(new_n583), .B2(new_n584), .C1(new_n698), .C2(new_n288), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n700), .ZN(new_n757));
  INV_X1    g0557(.A(new_n656), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n757), .A2(new_n531), .A3(new_n758), .A4(new_n713), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n737), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n564), .A2(new_n703), .A3(new_n581), .A4(new_n652), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n684), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n703), .B1(new_n700), .B2(new_n704), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT98), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n757), .A2(new_n765), .A3(new_n682), .A4(new_n687), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n755), .B1(new_n698), .B2(new_n288), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n586), .B(new_n687), .C1(new_n767), .C2(new_n580), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n653), .B1(G179), .B2(new_n612), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n595), .A2(new_n600), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n288), .ZN(new_n771));
  INV_X1    g0571(.A(new_n605), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n524), .A2(new_n530), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT98), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n764), .A2(new_n766), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(KEYINPUT29), .A3(new_n713), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT99), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n776), .A2(new_n779), .A3(KEYINPUT29), .A4(new_n713), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n705), .A2(new_n684), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n703), .B1(new_n700), .B2(new_n652), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n714), .B1(new_n784), .B2(new_n688), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT97), .B1(new_n785), .B2(KEYINPUT29), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n706), .A2(new_n713), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT97), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT29), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n760), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n736), .B1(new_n792), .B2(G1), .ZN(G364));
  AND2_X1   g0593(.A1(new_n210), .A2(G13), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G45), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n732), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n718), .B2(G330), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G330), .B2(new_n718), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  AOI21_X1  g0600(.A(new_n211), .B1(G20), .B2(new_n373), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n210), .A2(G179), .A3(G190), .A4(new_n311), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n297), .A2(new_n443), .A3(new_n311), .A4(G179), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT101), .Z(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n359), .B1(new_n802), .B2(new_n804), .C1(new_n807), .C2(new_n509), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G190), .A2(G200), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n545), .A2(new_n282), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G329), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n210), .A2(new_n282), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G190), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT33), .B(G317), .Z(new_n820));
  OAI22_X1  g0620(.A1(new_n814), .A2(new_n815), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n443), .A2(G200), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n210), .B1(new_n282), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n608), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n816), .A2(new_n809), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n816), .A2(new_n822), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n825), .B1(new_n826), .B2(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n817), .A2(new_n443), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(G326), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n808), .A2(new_n821), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n831), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n202), .A2(new_n834), .B1(new_n819), .B2(new_n224), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n810), .A2(KEYINPUT32), .A3(new_n350), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT32), .B1(new_n810), .B2(new_n350), .ZN(new_n837));
  INV_X1    g0637(.A(G58), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n836), .B(new_n837), .C1(new_n838), .C2(new_n829), .ZN(new_n839));
  INV_X1    g0639(.A(new_n805), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n275), .B1(new_n226), .B2(new_n840), .C1(new_n804), .C2(new_n231), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n824), .A2(G97), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n229), .B2(new_n826), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n835), .A2(new_n839), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n801), .B1(new_n833), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n359), .A2(new_n216), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n846), .A2(G355), .B1(new_n471), .B2(new_n216), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n247), .A2(new_n630), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n216), .A2(new_n325), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(G45), .B2(new_n207), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(G13), .A2(G33), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(G20), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n801), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n796), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n854), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n845), .B(new_n856), .C1(new_n718), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n800), .A2(new_n858), .ZN(G396));
  NOR2_X1   g0659(.A1(new_n410), .A2(new_n714), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n412), .B1(new_n407), .B2(new_n713), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n410), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n787), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n860), .B1(new_n410), .B2(new_n862), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n706), .A3(new_n713), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n760), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n797), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n804), .A2(new_n224), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n322), .B(new_n872), .C1(G58), .C2(new_n824), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n202), .B2(new_n807), .ZN(new_n874));
  INV_X1    g0674(.A(new_n826), .ZN(new_n875));
  INV_X1    g0675(.A(new_n829), .ZN(new_n876));
  AOI22_X1  g0676(.A1(G159), .A2(new_n875), .B1(new_n876), .B2(G143), .ZN(new_n877));
  INV_X1    g0677(.A(G137), .ZN(new_n878));
  INV_X1    g0678(.A(G150), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n877), .B1(new_n834), .B2(new_n878), .C1(new_n879), .C2(new_n819), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT34), .Z(new_n881));
  INV_X1    g0681(.A(new_n814), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n874), .B(new_n881), .C1(G132), .C2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n806), .A2(G107), .B1(G294), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n471), .B2(new_n826), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n275), .B1(new_n803), .B2(G87), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n842), .B(new_n886), .C1(new_n814), .C2(new_n827), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n802), .A2(new_n819), .B1(new_n834), .B2(new_n509), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n801), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n801), .A2(new_n852), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n796), .B1(new_n229), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n892), .C1(new_n853), .C2(new_n866), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n871), .A2(new_n893), .ZN(G384));
  NAND2_X1  g0694(.A1(new_n544), .A2(new_n550), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n897));
  INV_X1    g0697(.A(new_n211), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n898), .A4(new_n545), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n734), .A2(G77), .A3(new_n346), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n202), .A2(G68), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n255), .B(G13), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n470), .B1(new_n786), .B2(new_n790), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n781), .A2(new_n907), .A3(KEYINPUT105), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n677), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n778), .A2(new_n780), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(new_n912));
  AOI211_X1 g0712(.A(KEYINPUT97), .B(KEYINPUT29), .C1(new_n706), .C2(new_n713), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n678), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n910), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n663), .A2(new_n713), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n355), .A2(new_n288), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT78), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n353), .B1(new_n351), .B2(new_n352), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT16), .B1(new_n921), .B2(new_n344), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n369), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n712), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n387), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n370), .A2(new_n712), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n376), .A2(new_n927), .A3(new_n382), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n340), .A2(new_n375), .A3(new_n923), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n930), .A2(new_n382), .A3(new_n924), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n931), .B2(new_n927), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n926), .A2(new_n932), .A3(KEYINPUT38), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT104), .ZN(new_n938));
  INV_X1    g0738(.A(new_n928), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n387), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n376), .A2(new_n382), .A3(new_n928), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n929), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n938), .B1(new_n944), .B2(new_n934), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT39), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n387), .A2(new_n939), .B1(new_n942), .B2(new_n929), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n936), .B1(KEYINPUT38), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n917), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n860), .B1(new_n785), .B2(new_n863), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n431), .A2(new_n713), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n469), .B(new_n955), .C1(new_n671), .C2(new_n672), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n955), .B1(new_n461), .B2(new_n469), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n926), .A2(new_n932), .A3(KEYINPUT38), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n926), .B2(new_n932), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n953), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n666), .A2(new_n712), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n952), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n916), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n469), .B1(new_n671), .B2(new_n672), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n954), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n956), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n754), .A2(new_n759), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(new_n948), .A3(new_n971), .A4(new_n866), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT40), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n864), .B1(new_n969), .B2(new_n956), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT40), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n974), .A2(new_n937), .A3(new_n975), .A4(new_n971), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n470), .B1(new_n759), .B2(new_n754), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n737), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n967), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n255), .B2(new_n794), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n967), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n906), .B1(new_n982), .B2(new_n983), .ZN(G367));
  AOI21_X1  g0784(.A(new_n587), .B1(new_n564), .B2(new_n714), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n773), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n714), .B1(new_n986), .B2(new_n582), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n582), .A2(new_n713), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n728), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT42), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(KEYINPUT42), .A3(new_n728), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT106), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n628), .A2(new_n629), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n714), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(new_n684), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n704), .B2(new_n998), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(new_n994), .B2(KEYINPUT106), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT43), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT43), .A4(new_n995), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT107), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(KEYINPUT107), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n723), .A2(new_n989), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n795), .A2(G1), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n718), .A2(G330), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT111), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n726), .B2(new_n721), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1017), .B(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n728), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n792), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n729), .A2(new_n989), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n729), .B2(new_n989), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT110), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(KEYINPUT44), .C1(new_n729), .C2(new_n989), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(KEYINPUT44), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n729), .A2(new_n989), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT44), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(KEYINPUT110), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n724), .A2(new_n1028), .A3(new_n1030), .A4(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1030), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n723), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n792), .B1(new_n1022), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n731), .B(new_n1041), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n1016), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1010), .A2(new_n723), .A3(new_n989), .A4(new_n1011), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1014), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n801), .B(new_n854), .C1(new_n216), .C2(new_n643), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n242), .A2(new_n849), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n796), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n803), .A2(G97), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT114), .B(KEYINPUT46), .Z(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n840), .B2(new_n471), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n811), .A2(G317), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .A4(new_n322), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n806), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(G303), .C2(new_n876), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT113), .B(G311), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n608), .A2(new_n818), .B1(new_n831), .B2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n826), .A2(new_n802), .B1(new_n823), .B2(new_n231), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  NAND3_X1  g0859(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n823), .A2(new_n224), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G150), .B2(new_n876), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n202), .B2(new_n826), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n804), .A2(new_n229), .B1(new_n878), .B2(new_n810), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n359), .B(new_n1064), .C1(G58), .C2(new_n805), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n831), .A2(G143), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n350), .C2(new_n819), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1060), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT47), .Z(new_n1069));
  INV_X1    g0869(.A(new_n801), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1048), .B1(new_n857), .B2(new_n1001), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1045), .A2(new_n1071), .ZN(G387));
  OR2_X1    g0872(.A1(new_n239), .A2(new_n630), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n733), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1073), .A2(new_n849), .B1(new_n1074), .B2(new_n846), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n394), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1076), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n733), .B(new_n630), .C1(new_n224), .C2(new_n229), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT50), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n394), .B2(new_n202), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1075), .A2(new_n1081), .B1(G107), .B2(new_n215), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n796), .B1(new_n1082), .B2(new_n855), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n721), .B2(new_n857), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n325), .B1(new_n811), .B2(G326), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G303), .A2(new_n875), .B1(new_n876), .B2(G317), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n818), .A2(new_n1056), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n828), .C2(new_n834), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n824), .A2(G283), .B1(new_n805), .B2(new_n608), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT49), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1085), .B1(new_n471), .B2(new_n804), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n823), .A2(new_n396), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n826), .B2(new_n224), .C1(new_n202), .C2(new_n829), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1049), .B(new_n325), .C1(new_n229), .C2(new_n840), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G150), .B2(new_n811), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n818), .A2(new_n295), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n350), .C2(new_n834), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1095), .A2(new_n1096), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1084), .B1(new_n1104), .B2(new_n801), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT115), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1021), .B2(new_n1015), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1022), .A2(new_n731), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1021), .A2(new_n792), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(G393));
  OAI21_X1  g0910(.A(new_n855), .B1(new_n434), .B2(new_n215), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n250), .B2(new_n849), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT116), .ZN(new_n1113));
  INV_X1    g0913(.A(G294), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n826), .A2(new_n1114), .B1(new_n823), .B2(new_n471), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G107), .A2(new_n803), .B1(new_n811), .B2(G322), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1116), .B(new_n359), .C1(new_n802), .C2(new_n840), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G303), .C2(new_n818), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n831), .A2(G317), .B1(new_n876), .B2(G311), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT52), .Z(new_n1120));
  AOI22_X1  g0920(.A1(new_n831), .A2(G150), .B1(new_n876), .B2(G159), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT51), .Z(new_n1122));
  OAI22_X1  g0922(.A1(new_n826), .A2(new_n1076), .B1(new_n823), .B2(new_n229), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n811), .A2(G143), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n322), .B1(new_n805), .B2(G68), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n804), .C2(new_n226), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(G50), .C2(new_n818), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1118), .A2(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n797), .B(new_n1113), .C1(new_n1128), .C2(new_n1070), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n989), .B2(new_n857), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1038), .B2(new_n1016), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT118), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1021), .A2(new_n792), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n731), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n1139), .ZN(G390));
  INV_X1    g0940(.A(KEYINPUT39), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT104), .B1(new_n947), .B2(KEYINPUT38), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n962), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n948), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n853), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n807), .A2(new_n226), .B1(new_n471), .B2(new_n829), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G97), .B2(new_n875), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n882), .A2(G294), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n275), .B(new_n872), .C1(G77), .C2(new_n824), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G107), .A2(new_n818), .B1(new_n831), .B2(G283), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n805), .A2(G150), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n359), .B(new_n1153), .C1(G50), .C2(new_n803), .ZN(new_n1154));
  INV_X1    g0954(.A(G132), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1155), .A2(new_n829), .B1(new_n826), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G159), .B2(new_n824), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n882), .A2(G125), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n831), .B1(new_n818), .B2(G137), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1070), .B1(new_n1151), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n891), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n797), .B1(new_n295), .B2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1145), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n974), .A2(new_n760), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n917), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n867), .A2(new_n861), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n970), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1170), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n776), .A2(new_n713), .A3(new_n863), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n861), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1168), .B(new_n949), .C1(new_n1173), .C2(new_n970), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n970), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n917), .A3(new_n948), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n917), .B1(new_n953), .B2(new_n959), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n946), .A3(new_n951), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1179), .A3(new_n1166), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n1016), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1165), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n678), .A2(new_n760), .ZN(new_n1186));
  AND4_X1   g0986(.A1(new_n677), .A2(new_n915), .A3(new_n908), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT31), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n753), .B(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n759), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G330), .B(new_n866), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n959), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1166), .A2(new_n1192), .A3(new_n861), .A4(new_n1172), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1166), .A2(new_n1192), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(new_n953), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1187), .A2(new_n1195), .A3(new_n1175), .A4(new_n1180), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n909), .A2(new_n915), .A3(new_n1186), .A4(new_n1195), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1181), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n731), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1185), .A2(new_n1199), .ZN(G378));
  OAI21_X1  g1000(.A(new_n712), .B1(new_n303), .B2(new_n308), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n321), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1201), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n310), .B(new_n1203), .C1(new_n318), .C2(new_n320), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1206), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1202), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n970), .A2(new_n971), .A3(new_n866), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n962), .A2(KEYINPUT40), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1211), .A2(new_n1212), .B1(new_n972), .B2(KEYINPUT40), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1210), .B1(new_n1213), .B2(new_n737), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1210), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n977), .A2(new_n1215), .A3(G330), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1214), .A2(new_n965), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n965), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1210), .A2(new_n852), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n797), .B1(G50), .B2(new_n1163), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1061), .B1(new_n831), .B2(G116), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT120), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n803), .A2(G58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n322), .A2(new_n498), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G77), .B2(new_n805), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(new_n396), .C2(new_n826), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G107), .B2(new_n876), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n882), .A2(G283), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n818), .A2(G97), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1224), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT58), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G50), .B1(new_n271), .B2(new_n498), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1232), .A2(new_n1233), .B1(new_n1226), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n819), .A2(new_n1155), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n876), .A2(G128), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n875), .A2(G137), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n879), .B2(new_n823), .C1(new_n840), .C2(new_n1156), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1236), .B(new_n1240), .C1(G125), .C2(new_n831), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n803), .A2(G159), .ZN(new_n1244));
  AOI211_X1 g1044(.A(G33), .B(G41), .C1(new_n811), .C2(G124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1235), .B1(new_n1233), .B2(new_n1232), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(KEYINPUT121), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1070), .B1(new_n1248), .B2(KEYINPUT121), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1222), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1220), .A2(new_n1015), .B1(new_n1221), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT57), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT124), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n965), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n915), .A2(new_n677), .A3(new_n908), .A4(new_n1186), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT122), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT122), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n909), .A2(new_n1261), .A3(new_n915), .A4(new_n1186), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT123), .B1(new_n1263), .B2(new_n1196), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1260), .B(new_n1262), .C1(new_n1197), .C2(new_n1181), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT123), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1258), .B1(new_n1264), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n731), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1196), .A2(KEYINPUT123), .A3(new_n1260), .A4(new_n1262), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1272), .B2(new_n1220), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1252), .B1(new_n1269), .B2(new_n1273), .ZN(G375));
  NAND2_X1  g1074(.A1(new_n1195), .A2(new_n1015), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n882), .A2(G128), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n875), .A2(G150), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n325), .A3(new_n1225), .A4(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n806), .A2(G159), .B1(G50), .B2(new_n824), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n878), .B2(new_n829), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1155), .A2(new_n834), .B1(new_n819), .B2(new_n1156), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n806), .A2(G97), .B1(G107), .B2(new_n875), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n802), .B2(new_n829), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n814), .A2(new_n509), .B1(new_n819), .B2(new_n471), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n834), .A2(new_n1114), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1098), .B(new_n359), .C1(new_n229), .C2(new_n804), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n801), .B1(new_n1282), .B2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1289), .B(new_n797), .C1(G68), .C2(new_n1163), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(KEYINPUT125), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n970), .B2(new_n853), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1187), .A2(new_n1195), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1042), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1197), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1275), .B(new_n1292), .C1(new_n1293), .C2(new_n1295), .ZN(G381));
  OR4_X1    g1096(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1297), .A2(G387), .A3(G381), .ZN(new_n1298));
  INV_X1    g1098(.A(G378), .ZN(new_n1299));
  INV_X1    g1099(.A(G375), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(G407));
  INV_X1    g1101(.A(G343), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(G213), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(new_n1299), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G407), .A2(G213), .A3(new_n1305), .ZN(G409));
  OAI211_X1 g1106(.A(G378), .B(new_n1252), .C1(new_n1269), .C2(new_n1273), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1042), .B(new_n1219), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1251), .A2(new_n1221), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1016), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1299), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1307), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1303), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1197), .A2(KEYINPUT60), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1187), .B2(new_n1195), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1293), .A2(KEYINPUT60), .A3(new_n1197), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n731), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1275), .A2(new_n1292), .ZN(new_n1319));
  INV_X1    g1119(.A(G384), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(KEYINPUT126), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(KEYINPUT126), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1318), .B(new_n1321), .C1(KEYINPUT126), .C2(new_n1320), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1304), .A2(G2897), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1324), .A2(G2897), .A3(new_n1304), .A4(new_n1325), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1313), .A2(new_n1303), .A3(new_n1326), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  XOR2_X1   g1134(.A(G393), .B(G396), .Z(new_n1335));
  AOI21_X1  g1135(.A(G390), .B1(new_n1045), .B2(new_n1071), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1045), .A2(G390), .A3(new_n1071), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1335), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1045), .A2(G390), .A3(new_n1071), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1335), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1340), .A2(new_n1336), .A3(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1304), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(KEYINPUT63), .A3(new_n1326), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1331), .A2(new_n1334), .A3(new_n1343), .A4(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1347), .B1(new_n1344), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1332), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1344), .A2(KEYINPUT62), .A3(new_n1326), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1349), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1354), .B1(new_n1339), .B2(new_n1342), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1337), .A2(new_n1335), .A3(new_n1338), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1341), .B1(new_n1340), .B2(new_n1336), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1357), .A3(KEYINPUT127), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1346), .B1(new_n1353), .B2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1299), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1307), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1362), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1307), .A3(new_n1326), .ZN(new_n1364));
  AND3_X1   g1164(.A1(new_n1343), .A2(new_n1363), .A3(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1343), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(G402));
endmodule


