

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593;

  INV_X1 U322 ( .A(KEYINPUT112), .ZN(n393) );
  XNOR2_X1 U323 ( .A(n461), .B(KEYINPUT120), .ZN(n569) );
  XNOR2_X1 U324 ( .A(n584), .B(KEYINPUT41), .ZN(n558) );
  INV_X1 U325 ( .A(n558), .ZN(n568) );
  XOR2_X1 U326 ( .A(G29GAT), .B(G43GAT), .Z(n290) );
  XOR2_X1 U327 ( .A(KEYINPUT45), .B(n391), .Z(n291) );
  NAND2_X1 U328 ( .A1(n558), .A2(n553), .ZN(n349) );
  XNOR2_X1 U329 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U330 ( .A(n319), .B(n318), .ZN(n323) );
  XNOR2_X1 U331 ( .A(n394), .B(n393), .ZN(n395) );
  AND2_X1 U332 ( .A1(n396), .A2(n395), .ZN(n397) );
  NOR2_X1 U333 ( .A1(n425), .A2(n522), .ZN(n575) );
  XNOR2_X1 U334 ( .A(KEYINPUT48), .B(n397), .ZN(n552) );
  XOR2_X1 U335 ( .A(n366), .B(n365), .Z(n546) );
  XNOR2_X1 U336 ( .A(n465), .B(G190GAT), .ZN(n466) );
  XNOR2_X1 U337 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n442) );
  INV_X1 U339 ( .A(KEYINPUT54), .ZN(n400) );
  XOR2_X1 U340 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n293) );
  NAND2_X1 U341 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U343 ( .A(n294), .B(KEYINPUT94), .Z(n296) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .Z(n350) );
  XOR2_X1 U345 ( .A(G8GAT), .B(G183GAT), .Z(n378) );
  XNOR2_X1 U346 ( .A(n350), .B(n378), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n303) );
  INV_X1 U348 ( .A(G92GAT), .ZN(n297) );
  NAND2_X1 U349 ( .A1(G64GAT), .A2(n297), .ZN(n300) );
  INV_X1 U350 ( .A(G64GAT), .ZN(n298) );
  NAND2_X1 U351 ( .A1(n298), .A2(G92GAT), .ZN(n299) );
  NAND2_X1 U352 ( .A1(n300), .A2(n299), .ZN(n302) );
  XNOR2_X1 U353 ( .A(G176GAT), .B(G204GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n312) );
  XOR2_X1 U355 ( .A(n303), .B(n312), .Z(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n305) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n451) );
  XOR2_X1 U359 ( .A(KEYINPUT21), .B(G218GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(KEYINPUT87), .B(G211GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(G197GAT), .B(n308), .Z(n438) );
  XNOR2_X1 U363 ( .A(n451), .B(n438), .ZN(n309) );
  XOR2_X1 U364 ( .A(n310), .B(n309), .Z(n524) );
  INV_X1 U365 ( .A(n524), .ZN(n398) );
  XOR2_X1 U366 ( .A(G99GAT), .B(G85GAT), .Z(n351) );
  INV_X1 U367 ( .A(n312), .ZN(n311) );
  NAND2_X1 U368 ( .A1(n351), .A2(n311), .ZN(n315) );
  INV_X1 U369 ( .A(n351), .ZN(n313) );
  NAND2_X1 U370 ( .A1(n313), .A2(n312), .ZN(n314) );
  NAND2_X1 U371 ( .A1(n315), .A2(n314), .ZN(n319) );
  NAND2_X1 U372 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  INV_X1 U373 ( .A(KEYINPUT33), .ZN(n316) );
  XOR2_X1 U374 ( .A(G78GAT), .B(G148GAT), .Z(n321) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n428) );
  XNOR2_X1 U377 ( .A(n428), .B(KEYINPUT32), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U379 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n325) );
  XNOR2_X1 U380 ( .A(KEYINPUT31), .B(KEYINPUT75), .ZN(n324) );
  XOR2_X1 U381 ( .A(n325), .B(n324), .Z(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n329) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G71GAT), .ZN(n445) );
  XOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT13), .Z(n379) );
  XOR2_X1 U385 ( .A(n445), .B(n379), .Z(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n584) );
  XOR2_X1 U387 ( .A(G22GAT), .B(G141GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G50GAT), .B(G36GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G113GAT), .Z(n333) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G197GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U393 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n337) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U397 ( .A(KEYINPUT67), .B(n338), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U399 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n342) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n344), .B(n343), .Z(n348) );
  XNOR2_X1 U403 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n290), .B(n345), .ZN(n354) );
  XNOR2_X1 U405 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n346), .B(KEYINPUT70), .ZN(n375) );
  XNOR2_X1 U407 ( .A(n354), .B(n375), .ZN(n347) );
  XOR2_X1 U408 ( .A(n348), .B(n347), .Z(n553) );
  XNOR2_X1 U409 ( .A(n349), .B(KEYINPUT46), .ZN(n389) );
  XOR2_X1 U410 ( .A(n351), .B(n350), .Z(n353) );
  XOR2_X1 U411 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XOR2_X1 U412 ( .A(G134GAT), .B(KEYINPUT77), .Z(n415) );
  XNOR2_X1 U413 ( .A(n427), .B(n415), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U415 ( .A(G92GAT), .B(n354), .Z(n356) );
  NAND2_X1 U416 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U418 ( .A(n358), .B(n357), .Z(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n360) );
  XNOR2_X1 U420 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U422 ( .A(KEYINPUT65), .B(KEYINPUT64), .Z(n362) );
  XNOR2_X1 U423 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  INV_X1 U426 ( .A(n546), .ZN(n563) );
  XOR2_X1 U427 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n368) );
  XNOR2_X1 U428 ( .A(KEYINPUT79), .B(KEYINPUT81), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n387) );
  XOR2_X1 U430 ( .A(G64GAT), .B(G78GAT), .Z(n370) );
  XNOR2_X1 U431 ( .A(G71GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U433 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U434 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U436 ( .A(n374), .B(n373), .Z(n385) );
  XOR2_X1 U437 ( .A(n375), .B(KEYINPUT83), .Z(n377) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n383) );
  XOR2_X1 U440 ( .A(n379), .B(n378), .Z(n381) );
  XOR2_X1 U441 ( .A(G15GAT), .B(G127GAT), .Z(n446) );
  XOR2_X1 U442 ( .A(G22GAT), .B(G155GAT), .Z(n426) );
  XNOR2_X1 U443 ( .A(n446), .B(n426), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U447 ( .A(n387), .B(n386), .Z(n561) );
  NOR2_X1 U448 ( .A1(n563), .A2(n561), .ZN(n388) );
  AND2_X1 U449 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n390), .B(KEYINPUT47), .ZN(n396) );
  INV_X1 U451 ( .A(n553), .ZN(n576) );
  NAND2_X1 U452 ( .A1(n576), .A2(n584), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n546), .B(KEYINPUT36), .ZN(n591) );
  INV_X1 U454 ( .A(n561), .ZN(n588) );
  NOR2_X1 U455 ( .A1(n591), .A2(n588), .ZN(n391) );
  NOR2_X1 U456 ( .A1(n392), .A2(n291), .ZN(n394) );
  NOR2_X1 U457 ( .A1(n398), .A2(n552), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n425) );
  XOR2_X1 U459 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n402) );
  XNOR2_X1 U460 ( .A(G1GAT), .B(G120GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n404) );
  XNOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U465 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U466 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n408) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U469 ( .A(G57GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n419) );
  XOR2_X1 U471 ( .A(G148GAT), .B(G155GAT), .Z(n413) );
  XNOR2_X1 U472 ( .A(G127GAT), .B(G162GAT), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U474 ( .A(n414), .B(G85GAT), .Z(n417) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(n415), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n424) );
  XNOR2_X1 U478 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n420), .B(KEYINPUT84), .ZN(n447) );
  XOR2_X1 U480 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n422) );
  XNOR2_X1 U481 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n447), .B(n430), .ZN(n423) );
  XOR2_X1 U484 ( .A(n424), .B(n423), .Z(n480) );
  INV_X1 U485 ( .A(n480), .ZN(n522) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT22), .B(n430), .Z(n432) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U491 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n436) );
  XNOR2_X1 U493 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n476) );
  NAND2_X1 U497 ( .A1(n575), .A2(n476), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n460) );
  XOR2_X1 U499 ( .A(G190GAT), .B(G134GAT), .Z(n444) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G99GAT), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n459) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U503 ( .A(n448), .B(n447), .Z(n457) );
  XOR2_X1 U504 ( .A(KEYINPUT86), .B(G176GAT), .Z(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n455) );
  XOR2_X1 U507 ( .A(G183GAT), .B(n451), .Z(n453) );
  NAND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n536) );
  NAND2_X1 U513 ( .A1(n460), .A2(n536), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n569), .A2(n588), .ZN(n464) );
  INV_X1 U515 ( .A(G183GAT), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT122), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(G1350GAT) );
  NOR2_X1 U518 ( .A1(n569), .A2(n546), .ZN(n467) );
  INV_X1 U519 ( .A(KEYINPUT58), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n584), .A2(n553), .ZN(n498) );
  NOR2_X1 U521 ( .A1(n563), .A2(n588), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n468), .B(KEYINPUT16), .ZN(n484) );
  XNOR2_X1 U523 ( .A(n524), .B(KEYINPUT27), .ZN(n474) );
  NAND2_X1 U524 ( .A1(n474), .A2(n522), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT97), .ZN(n550) );
  XOR2_X1 U526 ( .A(n476), .B(KEYINPUT28), .Z(n530) );
  INV_X1 U527 ( .A(n530), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n550), .A2(n470), .ZN(n535) );
  NOR2_X1 U529 ( .A1(n536), .A2(n535), .ZN(n471) );
  XOR2_X1 U530 ( .A(KEYINPUT98), .B(n471), .Z(n483) );
  NOR2_X1 U531 ( .A1(n476), .A2(n536), .ZN(n472) );
  XOR2_X1 U532 ( .A(KEYINPUT26), .B(n472), .Z(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT99), .B(n473), .ZN(n574) );
  NAND2_X1 U534 ( .A1(n574), .A2(n474), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n536), .A2(n524), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT25), .B(n477), .Z(n478) );
  NAND2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n495) );
  NAND2_X1 U541 ( .A1(n484), .A2(n495), .ZN(n510) );
  NOR2_X1 U542 ( .A1(n498), .A2(n510), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT100), .B(n485), .ZN(n492) );
  NAND2_X1 U544 ( .A1(n492), .A2(n522), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT34), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  XOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT101), .Z(n489) );
  NAND2_X1 U548 ( .A1(n492), .A2(n524), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U551 ( .A1(n492), .A2(n536), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n492), .A2(n530), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT102), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n494), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n501) );
  NAND2_X1 U557 ( .A1(n588), .A2(n495), .ZN(n496) );
  NOR2_X1 U558 ( .A1(n591), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n497), .ZN(n521) );
  NOR2_X1 U560 ( .A1(n498), .A2(n521), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT38), .ZN(n507) );
  NAND2_X1 U562 ( .A1(n522), .A2(n507), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U564 ( .A(G29GAT), .B(n502), .Z(G1328GAT) );
  NAND2_X1 U565 ( .A1(n507), .A2(n524), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n505) );
  NAND2_X1 U568 ( .A1(n507), .A2(n536), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U570 ( .A(G43GAT), .B(n506), .Z(G1330GAT) );
  XOR2_X1 U571 ( .A(G50GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U572 ( .A1(n530), .A2(n507), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n512) );
  NAND2_X1 U575 ( .A1(n576), .A2(n558), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n510), .A2(n520), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n516), .A2(n522), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NAND2_X1 U580 ( .A1(n524), .A2(n516), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n536), .A2(n516), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n518) );
  NAND2_X1 U585 ( .A1(n516), .A2(n530), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n522), .A2(n531), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U592 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n536), .A2(n531), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(KEYINPUT110), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n533) );
  NAND2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n552), .A2(n535), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n545) );
  NOR2_X1 U604 ( .A1(n576), .A2(n545), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  NOR2_X1 U607 ( .A1(n568), .A2(n545), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U611 ( .A1(n588), .A2(n545), .ZN(n543) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n549), .Z(G1343GAT) );
  NAND2_X1 U618 ( .A1(n550), .A2(n574), .ZN(n551) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n553), .A2(n564), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT52), .B(n557), .Z(n560) );
  NAND2_X1 U626 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT118), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n576), .A2(n569), .ZN(n567) );
  XOR2_X1 U634 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n571) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n590) );
  NOR2_X1 U641 ( .A1(n576), .A2(n590), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT60), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n586) );
  NOR2_X1 U650 ( .A1(n584), .A2(n590), .ZN(n585) );
  XOR2_X1 U651 ( .A(n586), .B(n585), .Z(n587) );
  XNOR2_X1 U652 ( .A(KEYINPUT125), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

