//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1190, new_n1191;
  NOR2_X1   g000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g001(.A(G50), .ZN(new_n202));
  NAND2_X1  g002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  NOR2_X1   g005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g010(.A(G87), .ZN(new_n211));
  INV_X1    g011(.A(G250), .ZN(new_n212));
  INV_X1    g012(.A(G116), .ZN(new_n213));
  INV_X1    g013(.A(G270), .ZN(new_n214));
  OAI221_X1 g014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g015(.A(new_n215), .B1(G50), .B2(G226), .ZN(new_n216));
  INV_X1    g016(.A(G58), .ZN(new_n217));
  INV_X1    g017(.A(G232), .ZN(new_n218));
  INV_X1    g018(.A(G107), .ZN(new_n219));
  INV_X1    g019(.A(G264), .ZN(new_n220));
  OAI221_X1 g020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g021(.A(G68), .ZN(new_n222));
  INV_X1    g022(.A(G238), .ZN(new_n223));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g025(.A(new_n225), .B(KEYINPUT67), .Z(new_n226));
  XNOR2_X1  g026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  INV_X1    g027(.A(G20), .ZN(new_n228));
  NAND2_X1  g028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g032(.A1(G1), .A2(G13), .ZN(new_n233));
  OAI21_X1  g033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  NOR3_X1   g034(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g035(.A1(new_n209), .A2(G13), .ZN(new_n236));
  OAI211_X1 g036(.A(new_n236), .B(G250), .C1(G257), .C2(G264), .ZN(new_n237));
  XOR2_X1   g037(.A(new_n237), .B(KEYINPUT65), .Z(new_n238));
  XNOR2_X1  g038(.A(new_n238), .B(KEYINPUT0), .ZN(new_n239));
  NOR3_X1   g039(.A1(new_n227), .A2(new_n235), .A3(new_n239), .ZN(G361));
  XNOR2_X1  g040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g044(.A(G250), .B(G257), .Z(new_n245));
  XNOR2_X1  g045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g049(.A(new_n249), .B(new_n213), .ZN(new_n250));
  XOR2_X1   g050(.A(KEYINPUT68), .B(G107), .Z(new_n251));
  XNOR2_X1  g051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g052(.A(G68), .B(G77), .ZN(new_n253));
  XNOR2_X1  g053(.A(G50), .B(G58), .ZN(new_n254));
  XNOR2_X1  g054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g055(.A(new_n252), .B(new_n255), .Z(G351));
  NAND2_X1  g056(.A1(G33), .A2(G97), .ZN(new_n257));
  INV_X1    g057(.A(G1698), .ZN(new_n258));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  NAND2_X1  g059(.A1(new_n259), .A2(G232), .ZN(new_n260));
  NAND3_X1  g060(.A1(new_n259), .A2(G226), .A3(new_n258), .ZN(new_n261));
  AND2_X1   g061(.A1(new_n261), .A2(KEYINPUT73), .ZN(new_n262));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n258), .ZN(new_n263));
  INV_X1    g063(.A(G226), .ZN(new_n264));
  NOR3_X1   g064(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n264), .ZN(new_n265));
  OAI221_X1 g065(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n262), .C2(new_n265), .ZN(new_n266));
  INV_X1    g066(.A(G33), .ZN(new_n267));
  INV_X1    g067(.A(G41), .ZN(new_n268));
  NOR2_X1   g068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OR2_X1    g069(.A1(new_n269), .A2(new_n233), .ZN(new_n270));
  INV_X1    g070(.A(new_n270), .ZN(new_n271));
  INV_X1    g071(.A(G1), .ZN(new_n272));
  OAI21_X1  g072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  AND2_X1   g073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g074(.A1(new_n266), .A2(new_n271), .B1(G238), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g075(.A1(new_n272), .A2(G274), .ZN(new_n276));
  OR2_X1    g076(.A1(KEYINPUT69), .A2(G41), .ZN(new_n277));
  NAND2_X1  g077(.A1(KEYINPUT69), .A2(G41), .ZN(new_n278));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g079(.A(G45), .ZN(new_n280));
  AOI21_X1  g080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g083(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n284));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n285));
  AOI21_X1  g085(.A(new_n285), .B1(new_n275), .B2(new_n282), .ZN(new_n286));
  OAI21_X1  g086(.A(G169), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g088(.A(new_n284), .ZN(new_n289));
  INV_X1    g089(.A(new_n286), .ZN(new_n290));
  NAND3_X1  g090(.A1(new_n289), .A2(G179), .A3(new_n290), .ZN(new_n291));
  INV_X1    g091(.A(KEYINPUT14), .ZN(new_n292));
  OAI211_X1 g092(.A(new_n292), .B(G169), .C1(new_n284), .C2(new_n286), .ZN(new_n293));
  NAND3_X1  g093(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g094(.A1(G20), .A2(G33), .ZN(new_n295));
  NAND2_X1  g095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NAND2_X1  g096(.A1(new_n232), .A2(G33), .ZN(new_n297));
  INV_X1    g097(.A(G77), .ZN(new_n298));
  OAI221_X1 g098(.A(new_n296), .B1(new_n228), .B2(G68), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  AND2_X1   g100(.A1(new_n300), .A2(new_n233), .ZN(new_n301));
  INV_X1    g101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g103(.A(new_n303), .B(KEYINPUT11), .Z(new_n304));
  AOI21_X1  g104(.A(new_n302), .B1(new_n272), .B2(G20), .ZN(new_n305));
  INV_X1    g105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n222), .ZN(new_n307));
  NAND3_X1  g107(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n308));
  INV_X1    g108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n222), .ZN(new_n310));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n311));
  XNOR2_X1  g111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NOR3_X1   g112(.A1(new_n304), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  INV_X1    g113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g115(.A1(new_n203), .A2(G20), .ZN(new_n316));
  INV_X1    g116(.A(G150), .ZN(new_n317));
  INV_X1    g117(.A(new_n295), .ZN(new_n318));
  XOR2_X1   g118(.A(KEYINPUT8), .B(G58), .Z(new_n319));
  INV_X1    g119(.A(new_n319), .ZN(new_n320));
  OAI221_X1 g120(.A(new_n316), .B1(new_n317), .B2(new_n318), .C1(new_n320), .C2(new_n297), .ZN(new_n321));
  AOI22_X1  g121(.A1(new_n321), .A2(new_n302), .B1(new_n202), .B2(new_n309), .ZN(new_n322));
  OAI21_X1  g122(.A(new_n322), .B1(new_n202), .B2(new_n306), .ZN(new_n323));
  XNOR2_X1  g123(.A(new_n323), .B(KEYINPUT9), .ZN(new_n324));
  INV_X1    g124(.A(new_n259), .ZN(new_n325));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n298), .ZN(new_n326));
  MUX2_X1   g126(.A(G222), .B(G223), .S(G1698), .Z(new_n327));
  OAI211_X1 g127(.A(new_n271), .B(new_n326), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g128(.A1(new_n270), .A2(new_n273), .ZN(new_n329));
  OAI211_X1 g129(.A(new_n328), .B(new_n282), .C1(new_n264), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  INV_X1    g131(.A(G190), .ZN(new_n332));
  OAI211_X1 g132(.A(new_n324), .B(new_n331), .C1(new_n332), .C2(new_n330), .ZN(new_n333));
  XNOR2_X1  g133(.A(new_n333), .B(KEYINPUT10), .ZN(new_n334));
  OR3_X1    g134(.A1(new_n330), .A2(KEYINPUT70), .A3(G179), .ZN(new_n335));
  INV_X1    g135(.A(G169), .ZN(new_n336));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g137(.A(KEYINPUT70), .B1(new_n330), .B2(G179), .ZN(new_n338));
  NAND4_X1  g138(.A1(new_n335), .A2(new_n323), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  AND2_X1   g139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g140(.A1(new_n289), .A2(new_n290), .ZN(new_n341));
  AOI21_X1  g141(.A(new_n314), .B1(new_n341), .B2(G200), .ZN(new_n342));
  OAI21_X1  g142(.A(new_n342), .B1(new_n332), .B2(new_n341), .ZN(new_n343));
  XNOR2_X1  g143(.A(KEYINPUT66), .B(G20), .ZN(new_n344));
  AOI22_X1  g144(.A1(new_n319), .A2(new_n295), .B1(new_n344), .B2(G77), .ZN(new_n345));
  XOR2_X1   g145(.A(new_n345), .B(KEYINPUT72), .Z(new_n346));
  XOR2_X1   g146(.A(KEYINPUT15), .B(G87), .Z(new_n347));
  INV_X1    g147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g148(.A(new_n346), .B1(new_n297), .B2(new_n348), .ZN(new_n349));
  AOI22_X1  g149(.A1(new_n349), .A2(new_n302), .B1(new_n298), .B2(new_n309), .ZN(new_n350));
  OAI21_X1  g150(.A(new_n350), .B1(new_n298), .B2(new_n306), .ZN(new_n351));
  AOI21_X1  g151(.A(new_n281), .B1(new_n274), .B2(G244), .ZN(new_n352));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n353));
  OR2_X1    g153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g154(.A1(new_n259), .A2(G1698), .ZN(new_n355));
  OAI22_X1  g155(.A1(new_n355), .A2(new_n223), .B1(new_n219), .B2(new_n259), .ZN(new_n356));
  NOR2_X1   g156(.A1(new_n260), .A2(G1698), .ZN(new_n357));
  OAI21_X1  g157(.A(new_n271), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g158(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g160(.A(new_n351), .B1(G200), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g161(.A(new_n361), .B1(new_n332), .B2(new_n360), .ZN(new_n362));
  AND4_X1   g162(.A1(new_n315), .A2(new_n340), .A3(new_n343), .A4(new_n362), .ZN(new_n363));
  XNOR2_X1  g163(.A(G58), .B(G68), .ZN(new_n364));
  AOI22_X1  g164(.A1(new_n364), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n365));
  NAND2_X1  g165(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g167(.A1(new_n367), .A2(G33), .ZN(new_n368));
  AOI22_X1  g168(.A1(new_n229), .A2(new_n231), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g169(.A(KEYINPUT74), .B1(new_n369), .B2(KEYINPUT7), .ZN(new_n370));
  AOI21_X1  g170(.A(G20), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g171(.A1(new_n371), .A2(KEYINPUT7), .ZN(new_n372));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n373));
  INV_X1    g173(.A(KEYINPUT7), .ZN(new_n374));
  OAI211_X1 g174(.A(new_n373), .B(new_n374), .C1(new_n344), .C2(new_n259), .ZN(new_n375));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT75), .A3(G68), .ZN(new_n377));
  AOI21_X1  g177(.A(KEYINPUT75), .B1(new_n376), .B2(G68), .ZN(new_n378));
  OAI211_X1 g178(.A(KEYINPUT16), .B(new_n365), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NOR2_X1   g179(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n380));
  NOR2_X1   g180(.A1(new_n367), .A2(G33), .ZN(new_n381));
  AOI21_X1  g181(.A(new_n380), .B1(KEYINPUT77), .B2(new_n381), .ZN(new_n382));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g184(.A(new_n344), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n386));
  OAI21_X1  g186(.A(new_n386), .B1(new_n371), .B2(KEYINPUT7), .ZN(new_n387));
  OAI211_X1 g187(.A(KEYINPUT76), .B(new_n374), .C1(new_n259), .C2(G20), .ZN(new_n388));
  AOI22_X1  g188(.A1(new_n385), .A2(KEYINPUT7), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g189(.A(new_n365), .B1(new_n389), .B2(new_n222), .ZN(new_n390));
  INV_X1    g190(.A(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g191(.A(new_n301), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g192(.A1(new_n379), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g193(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  NOR2_X1   g194(.A1(new_n319), .A2(new_n309), .ZN(new_n395));
  AOI21_X1  g195(.A(new_n395), .B1(new_n306), .B2(new_n319), .ZN(new_n396));
  INV_X1    g196(.A(new_n396), .ZN(new_n397));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n398));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n398), .A3(new_n392), .ZN(new_n399));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g200(.A(new_n282), .B1(new_n329), .B2(new_n218), .ZN(new_n401));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n402));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g203(.A(new_n282), .B(KEYINPUT79), .C1(new_n329), .C2(new_n218), .ZN(new_n404));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g205(.A1(new_n264), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g206(.A(new_n259), .B(new_n406), .C1(G223), .C2(G1698), .ZN(new_n407));
  NAND2_X1  g207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g208(.A(new_n270), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g210(.A(G179), .ZN(new_n411));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g212(.A(new_n336), .B1(new_n401), .B2(new_n409), .ZN(new_n413));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g214(.A(new_n414), .ZN(new_n415));
  AND3_X1   g215(.A1(new_n400), .A2(KEYINPUT18), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g216(.A(KEYINPUT18), .B1(new_n400), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n332), .ZN(new_n419));
  INV_X1    g219(.A(G200), .ZN(new_n420));
  OAI21_X1  g220(.A(new_n420), .B1(new_n401), .B2(new_n409), .ZN(new_n421));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g222(.A1(new_n394), .A2(new_n422), .A3(new_n397), .A4(new_n399), .ZN(new_n423));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n424));
  XNOR2_X1  g224(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NOR2_X1   g225(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g226(.A1(new_n360), .A2(new_n336), .ZN(new_n427));
  OAI211_X1 g227(.A(new_n351), .B(new_n427), .C1(G179), .C2(new_n360), .ZN(new_n428));
  AND3_X1   g228(.A1(new_n363), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g230(.A1(new_n272), .A2(G33), .ZN(new_n431));
  NAND3_X1  g231(.A1(new_n301), .A2(new_n308), .A3(new_n431), .ZN(new_n432));
  INV_X1    g232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g233(.A1(new_n433), .A2(G116), .ZN(new_n434));
  NAND2_X1  g234(.A1(G33), .A2(G283), .ZN(new_n435));
  INV_X1    g235(.A(G97), .ZN(new_n436));
  OAI211_X1 g236(.A(new_n232), .B(new_n435), .C1(G33), .C2(new_n436), .ZN(new_n437));
  OAI211_X1 g237(.A(new_n437), .B(new_n302), .C1(new_n228), .C2(G116), .ZN(new_n438));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n439));
  AND2_X1   g239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g240(.A1(new_n438), .A2(new_n439), .ZN(new_n441));
  OAI221_X1 g241(.A(new_n434), .B1(G116), .B2(new_n308), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g242(.A(new_n442), .ZN(new_n443));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n444));
  NAND3_X1  g244(.A1(new_n277), .A2(new_n444), .A3(new_n278), .ZN(new_n445));
  NOR2_X1   g245(.A1(new_n280), .A2(G1), .ZN(new_n446));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n448));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g249(.A1(new_n445), .A2(KEYINPUT80), .A3(new_n446), .ZN(new_n450));
  AND2_X1   g250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g251(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n452));
  NAND4_X1  g252(.A1(new_n451), .A2(G274), .A3(new_n270), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g253(.A1(new_n325), .A2(G303), .ZN(new_n454));
  INV_X1    g254(.A(G257), .ZN(new_n455));
  OAI221_X1 g255(.A(new_n454), .B1(new_n263), .B2(new_n455), .C1(new_n220), .C2(new_n355), .ZN(new_n456));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n271), .ZN(new_n457));
  NAND3_X1  g257(.A1(new_n449), .A2(new_n452), .A3(new_n450), .ZN(new_n458));
  NAND3_X1  g258(.A1(new_n458), .A2(G270), .A3(new_n270), .ZN(new_n459));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  OAI21_X1  g261(.A(KEYINPUT21), .B1(new_n443), .B2(new_n461), .ZN(new_n462));
  INV_X1    g262(.A(KEYINPUT21), .ZN(new_n463));
  NAND4_X1  g263(.A1(new_n442), .A2(new_n460), .A3(new_n463), .A4(G169), .ZN(new_n464));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g265(.A1(new_n443), .A2(new_n411), .A3(new_n460), .ZN(new_n466));
  INV_X1    g266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g267(.A1(new_n460), .A2(G200), .ZN(new_n468));
  OAI211_X1 g268(.A(new_n443), .B(new_n468), .C1(new_n332), .C2(new_n460), .ZN(new_n469));
  AND3_X1   g269(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n471));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n472));
  NOR2_X1   g272(.A1(new_n472), .A2(KEYINPUT24), .ZN(new_n473));
  NAND3_X1  g273(.A1(new_n232), .A2(new_n259), .A3(G87), .ZN(new_n474));
  NAND2_X1  g274(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n475));
  INV_X1    g275(.A(KEYINPUT22), .ZN(new_n476));
  NAND4_X1  g276(.A1(new_n232), .A2(new_n259), .A3(new_n476), .A4(G87), .ZN(new_n477));
  AND2_X1   g277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n479));
  NAND4_X1  g279(.A1(new_n229), .A2(new_n231), .A3(new_n479), .A4(new_n219), .ZN(new_n480));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g282(.A1(new_n344), .A2(KEYINPUT83), .A3(new_n479), .A4(new_n219), .ZN(new_n483));
  OAI21_X1  g283(.A(KEYINPUT23), .B1(new_n228), .B2(G107), .ZN(new_n484));
  INV_X1    g284(.A(KEYINPUT82), .ZN(new_n485));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g286(.A(KEYINPUT82), .B(KEYINPUT23), .C1(new_n228), .C2(G107), .ZN(new_n487));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g288(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n489));
  NAND4_X1  g289(.A1(new_n482), .A2(new_n483), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  OAI21_X1  g290(.A(new_n473), .B1(new_n478), .B2(new_n490), .ZN(new_n491));
  AND4_X1   g291(.A1(new_n483), .A2(new_n482), .A3(new_n488), .A4(new_n489), .ZN(new_n492));
  INV_X1    g292(.A(new_n473), .ZN(new_n493));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n477), .ZN(new_n494));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g295(.A1(new_n491), .A2(new_n495), .B1(new_n472), .B2(KEYINPUT24), .ZN(new_n496));
  OAI21_X1  g296(.A(new_n471), .B1(new_n496), .B2(new_n301), .ZN(new_n497));
  NAND2_X1  g297(.A1(new_n472), .A2(KEYINPUT24), .ZN(new_n498));
  NOR3_X1   g298(.A1(new_n478), .A2(new_n473), .A3(new_n490), .ZN(new_n499));
  AOI21_X1  g299(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n500));
  OAI21_X1  g300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n302), .ZN(new_n502));
  OAI21_X1  g302(.A(KEYINPUT87), .B1(new_n308), .B2(G107), .ZN(new_n503));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n504));
  OR2_X1    g304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g305(.A1(new_n433), .A2(G107), .ZN(new_n506));
  NAND4_X1  g306(.A1(new_n497), .A2(new_n502), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  OR3_X1    g307(.A1(new_n308), .A2(KEYINPUT87), .A3(G107), .ZN(new_n508));
  AND3_X1   g308(.A1(new_n508), .A2(new_n503), .A3(new_n504), .ZN(new_n509));
  NOR2_X1   g309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g310(.A1(G33), .A2(G294), .ZN(new_n511));
  OAI221_X1 g311(.A(new_n511), .B1(new_n263), .B2(new_n212), .C1(new_n455), .C2(new_n355), .ZN(new_n512));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n271), .ZN(new_n513));
  AND2_X1   g313(.A1(new_n453), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g314(.A1(new_n458), .A2(G264), .A3(new_n270), .ZN(new_n515));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g317(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  AND3_X1   g318(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g319(.A1(new_n514), .A2(new_n515), .ZN(new_n520));
  OAI22_X1  g320(.A1(new_n519), .A2(G200), .B1(G190), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g321(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g322(.A1(new_n433), .A2(G97), .ZN(new_n523));
  NAND2_X1  g323(.A1(new_n309), .A2(new_n436), .ZN(new_n524));
  NAND2_X1  g324(.A1(new_n387), .A2(new_n388), .ZN(new_n525));
  INV_X1    g325(.A(new_n384), .ZN(new_n526));
  OAI21_X1  g326(.A(new_n368), .B1(new_n366), .B2(new_n383), .ZN(new_n527));
  OAI211_X1 g327(.A(KEYINPUT7), .B(new_n232), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AOI21_X1  g328(.A(new_n219), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g329(.A1(new_n318), .A2(new_n298), .ZN(new_n530));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n531));
  NOR2_X1   g331(.A1(new_n436), .A2(new_n219), .ZN(new_n532));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n206), .ZN(new_n533));
  NAND3_X1  g333(.A1(new_n219), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  AND2_X1   g334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n232), .ZN(new_n536));
  NOR3_X1   g336(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g337(.A(new_n523), .B(new_n524), .C1(new_n537), .C2(new_n301), .ZN(new_n538));
  INV_X1    g338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g339(.A1(new_n458), .A2(G257), .A3(new_n270), .ZN(new_n540));
  NAND3_X1  g340(.A1(new_n259), .A2(G244), .A3(new_n258), .ZN(new_n541));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g343(.A(new_n543), .B1(new_n212), .B2(new_n355), .ZN(new_n544));
  OAI21_X1  g344(.A(new_n435), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g345(.A(new_n271), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g346(.A1(new_n453), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  INV_X1    g348(.A(new_n547), .ZN(new_n549));
  NAND2_X1  g349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  NAND3_X1  g350(.A1(new_n539), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n336), .ZN(new_n552));
  NAND4_X1  g352(.A1(new_n453), .A2(new_n411), .A3(new_n546), .A4(new_n540), .ZN(new_n553));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g354(.A1(new_n347), .A2(new_n308), .ZN(new_n555));
  NOR2_X1   g355(.A1(new_n432), .A2(new_n211), .ZN(new_n556));
  NAND3_X1  g356(.A1(new_n232), .A2(new_n259), .A3(G68), .ZN(new_n557));
  AND3_X1   g357(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n558));
  OAI22_X1  g358(.A1(new_n344), .A2(new_n558), .B1(G87), .B2(new_n207), .ZN(new_n559));
  NOR3_X1   g359(.A1(new_n344), .A2(new_n267), .A3(new_n436), .ZN(new_n560));
  OAI211_X1 g360(.A(new_n557), .B(new_n559), .C1(new_n560), .C2(KEYINPUT19), .ZN(new_n561));
  AOI211_X1 g361(.A(new_n555), .B(new_n556), .C1(new_n561), .C2(new_n302), .ZN(new_n562));
  NAND4_X1  g362(.A1(new_n366), .A2(new_n368), .A3(G244), .A4(G1698), .ZN(new_n563));
  NAND2_X1  g363(.A1(new_n563), .A2(KEYINPUT81), .ZN(new_n564));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n565));
  NAND4_X1  g365(.A1(new_n259), .A2(new_n565), .A3(G244), .A4(G1698), .ZN(new_n566));
  NAND2_X1  g366(.A1(G33), .A2(G116), .ZN(new_n567));
  NAND3_X1  g367(.A1(new_n259), .A2(G238), .A3(new_n258), .ZN(new_n568));
  NAND4_X1  g368(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n271), .ZN(new_n570));
  NOR2_X1   g370(.A1(new_n276), .A2(new_n280), .ZN(new_n571));
  INV_X1    g371(.A(new_n571), .ZN(new_n572));
  OAI221_X1 g372(.A(G250), .B1(G1), .B2(new_n280), .C1(new_n269), .C2(new_n233), .ZN(new_n573));
  NAND4_X1  g373(.A1(new_n570), .A2(G190), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  INV_X1    g374(.A(new_n573), .ZN(new_n575));
  AOI211_X1 g375(.A(new_n571), .B(new_n575), .C1(new_n569), .C2(new_n271), .ZN(new_n576));
  OAI211_X1 g376(.A(new_n562), .B(new_n574), .C1(new_n576), .C2(new_n420), .ZN(new_n577));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n302), .ZN(new_n578));
  INV_X1    g378(.A(new_n555), .ZN(new_n579));
  NAND2_X1  g379(.A1(new_n433), .A2(new_n347), .ZN(new_n580));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g381(.A1(new_n570), .A2(new_n411), .A3(new_n572), .A4(new_n573), .ZN(new_n582));
  OAI211_X1 g382(.A(new_n581), .B(new_n582), .C1(new_n576), .C2(G169), .ZN(new_n583));
  AND2_X1   g383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g384(.A1(new_n551), .A2(new_n554), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g385(.A1(new_n520), .A2(G169), .ZN(new_n586));
  NAND3_X1  g386(.A1(new_n514), .A2(new_n518), .A3(new_n517), .ZN(new_n587));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n411), .ZN(new_n588));
  OAI21_X1  g388(.A(new_n588), .B1(new_n507), .B2(new_n509), .ZN(new_n589));
  NAND4_X1  g389(.A1(new_n470), .A2(new_n522), .A3(new_n585), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g390(.A1(new_n430), .A2(new_n590), .ZN(G372));
  INV_X1    g391(.A(new_n339), .ZN(new_n592));
  INV_X1    g392(.A(new_n418), .ZN(new_n593));
  NAND2_X1  g393(.A1(new_n315), .A2(new_n428), .ZN(new_n594));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n343), .ZN(new_n595));
  OAI21_X1  g395(.A(new_n593), .B1(new_n595), .B2(new_n425), .ZN(new_n596));
  AOI21_X1  g396(.A(new_n592), .B1(new_n596), .B2(new_n334), .ZN(new_n597));
  AOI21_X1  g397(.A(new_n466), .B1(new_n462), .B2(new_n464), .ZN(new_n598));
  NAND2_X1  g398(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n585), .A3(new_n522), .ZN(new_n600));
  NAND2_X1  g400(.A1(new_n600), .A2(KEYINPUT89), .ZN(new_n601));
  INV_X1    g401(.A(KEYINPUT26), .ZN(new_n602));
  NAND2_X1  g402(.A1(new_n577), .A2(new_n583), .ZN(new_n603));
  OAI21_X1  g403(.A(new_n602), .B1(new_n554), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g404(.A1(new_n535), .A2(new_n232), .ZN(new_n605));
  INV_X1    g405(.A(new_n530), .ZN(new_n606));
  OAI211_X1 g406(.A(new_n605), .B(new_n606), .C1(new_n389), .C2(new_n219), .ZN(new_n607));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n302), .B1(new_n436), .B2(new_n309), .ZN(new_n608));
  AOI22_X1  g408(.A1(new_n608), .A2(new_n523), .B1(new_n547), .B2(new_n336), .ZN(new_n609));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n584), .A3(KEYINPUT26), .A4(new_n553), .ZN(new_n610));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n583), .ZN(new_n612));
  NAND2_X1  g412(.A1(new_n612), .A2(KEYINPUT90), .ZN(new_n613));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n614));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n614), .A3(new_n583), .ZN(new_n615));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g416(.A(KEYINPUT89), .ZN(new_n617));
  NAND4_X1  g417(.A1(new_n599), .A2(new_n585), .A3(new_n522), .A4(new_n617), .ZN(new_n618));
  AND3_X1   g418(.A1(new_n601), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g419(.A(new_n597), .B1(new_n430), .B2(new_n619), .ZN(G369));
  NAND2_X1  g420(.A1(new_n522), .A2(new_n589), .ZN(new_n621));
  INV_X1    g421(.A(new_n621), .ZN(new_n622));
  INV_X1    g422(.A(G13), .ZN(new_n623));
  NOR2_X1   g423(.A1(new_n344), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n272), .ZN(new_n625));
  OR2_X1    g425(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n626));
  NAND2_X1  g426(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n627));
  NAND3_X1  g427(.A1(new_n626), .A2(G213), .A3(new_n627), .ZN(new_n628));
  INV_X1    g428(.A(G343), .ZN(new_n629));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g431(.A(new_n622), .B1(new_n510), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g432(.A(new_n632), .B1(new_n589), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g433(.A1(new_n598), .A2(new_n630), .ZN(new_n634));
  OR2_X1    g434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g435(.A1(new_n443), .A2(new_n631), .ZN(new_n636));
  INV_X1    g436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g437(.A1(new_n470), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g438(.A1(new_n598), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g442(.A1(new_n622), .A2(new_n634), .ZN(new_n643));
  AND2_X1   g443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g444(.A(new_n589), .ZN(new_n645));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n631), .ZN(new_n646));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n646), .ZN(G399));
  INV_X1    g447(.A(new_n279), .ZN(new_n648));
  INV_X1    g448(.A(new_n236), .ZN(new_n649));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g451(.A1(new_n206), .A2(new_n211), .A3(new_n213), .ZN(new_n652));
  XNOR2_X1  g452(.A(new_n652), .B(KEYINPUT91), .ZN(new_n653));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n653), .A3(G1), .ZN(new_n654));
  OAI21_X1  g454(.A(new_n654), .B1(new_n234), .B2(new_n651), .ZN(new_n655));
  XNOR2_X1  g455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  NOR2_X1   g456(.A1(new_n619), .A2(new_n630), .ZN(new_n657));
  INV_X1    g457(.A(KEYINPUT92), .ZN(new_n658));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g459(.A(KEYINPUT29), .ZN(new_n660));
  INV_X1    g460(.A(new_n612), .ZN(new_n661));
  AOI21_X1  g461(.A(new_n630), .B1(new_n600), .B2(new_n661), .ZN(new_n662));
  NOR3_X1   g462(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g463(.A(new_n657), .ZN(new_n664));
  AOI21_X1  g464(.A(KEYINPUT29), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  NOR2_X1   g465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g466(.A1(new_n587), .A2(new_n411), .ZN(new_n667));
  NAND2_X1  g467(.A1(new_n546), .A2(new_n540), .ZN(new_n668));
  NOR2_X1   g468(.A1(new_n460), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n576), .A3(new_n669), .ZN(new_n670));
  INV_X1    g470(.A(KEYINPUT30), .ZN(new_n671));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g472(.A1(new_n667), .A2(KEYINPUT30), .A3(new_n576), .A4(new_n669), .ZN(new_n673));
  NAND4_X1  g473(.A1(new_n587), .A2(new_n411), .A3(new_n460), .A4(new_n547), .ZN(new_n674));
  OAI211_X1 g474(.A(new_n672), .B(new_n673), .C1(new_n576), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n630), .ZN(new_n676));
  OR2_X1    g476(.A1(new_n676), .A2(KEYINPUT31), .ZN(new_n677));
  OAI211_X1 g477(.A(new_n676), .B(KEYINPUT31), .C1(new_n590), .C2(new_n630), .ZN(new_n678));
  AND2_X1   g478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n680), .ZN(new_n681));
  INV_X1    g481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g482(.A(new_n656), .B1(new_n682), .B2(G1), .ZN(G364));
  NOR2_X1   g483(.A1(new_n640), .A2(G330), .ZN(new_n684));
  AOI21_X1  g484(.A(new_n272), .B1(new_n624), .B2(G45), .ZN(new_n685));
  INV_X1    g485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n650), .ZN(new_n687));
  OR3_X1    g487(.A1(new_n641), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  INV_X1    g488(.A(new_n687), .ZN(new_n689));
  NOR2_X1   g489(.A1(new_n232), .A2(G190), .ZN(new_n690));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n411), .A3(new_n420), .ZN(new_n691));
  OR2_X1    g491(.A1(new_n691), .A2(KEYINPUT94), .ZN(new_n692));
  NAND2_X1  g492(.A1(new_n691), .A2(KEYINPUT94), .ZN(new_n693));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g495(.A1(new_n344), .A2(G179), .A3(G190), .ZN(new_n696));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n420), .ZN(new_n697));
  AOI22_X1  g497(.A1(new_n695), .A2(G329), .B1(G326), .B2(new_n697), .ZN(new_n698));
  INV_X1    g498(.A(G294), .ZN(new_n699));
  NOR3_X1   g499(.A1(new_n332), .A2(G179), .A3(G200), .ZN(new_n700));
  NOR2_X1   g500(.A1(new_n232), .A2(new_n700), .ZN(new_n701));
  INV_X1    g501(.A(G311), .ZN(new_n702));
  NAND2_X1  g502(.A1(new_n690), .A2(G179), .ZN(new_n703));
  NOR2_X1   g503(.A1(new_n703), .A2(G200), .ZN(new_n704));
  INV_X1    g504(.A(new_n704), .ZN(new_n705));
  OAI221_X1 g505(.A(new_n698), .B1(new_n699), .B2(new_n701), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  NOR2_X1   g506(.A1(new_n703), .A2(new_n420), .ZN(new_n707));
  XNOR2_X1  g507(.A(KEYINPUT33), .B(G317), .ZN(new_n708));
  AOI21_X1  g508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g509(.A1(new_n420), .A2(G179), .ZN(new_n710));
  NAND3_X1  g510(.A1(new_n710), .A2(G20), .A3(G190), .ZN(new_n711));
  OR2_X1    g511(.A1(new_n711), .A2(KEYINPUT96), .ZN(new_n712));
  NAND2_X1  g512(.A1(new_n711), .A2(KEYINPUT96), .ZN(new_n713));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g515(.A1(new_n715), .A2(G303), .ZN(new_n716));
  NOR2_X1   g516(.A1(new_n696), .A2(G200), .ZN(new_n717));
  NAND2_X1  g517(.A1(new_n717), .A2(G322), .ZN(new_n718));
  NAND2_X1  g518(.A1(new_n690), .A2(new_n710), .ZN(new_n719));
  INV_X1    g519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g520(.A(new_n259), .B1(new_n720), .B2(G283), .ZN(new_n721));
  NAND4_X1  g521(.A1(new_n709), .A2(new_n716), .A3(new_n718), .A4(new_n721), .ZN(new_n722));
  INV_X1    g522(.A(new_n697), .ZN(new_n723));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n202), .ZN(new_n724));
  INV_X1    g524(.A(new_n707), .ZN(new_n725));
  OAI22_X1  g525(.A1(new_n222), .A2(new_n725), .B1(new_n705), .B2(new_n298), .ZN(new_n726));
  AOI211_X1 g526(.A(new_n724), .B(new_n726), .C1(G58), .C2(new_n717), .ZN(new_n727));
  INV_X1    g527(.A(G159), .ZN(new_n728));
  NOR2_X1   g528(.A1(new_n694), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g529(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n730));
  XNOR2_X1  g530(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g531(.A1(new_n720), .A2(G107), .ZN(new_n732));
  NAND3_X1  g532(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI221_X1 g533(.A(new_n259), .B1(new_n436), .B2(new_n701), .C1(new_n714), .C2(new_n211), .ZN(new_n734));
  OAI21_X1  g534(.A(new_n722), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g535(.A(KEYINPUT93), .B(G169), .ZN(new_n736));
  AOI21_X1  g536(.A(new_n233), .B1(new_n736), .B2(G20), .ZN(new_n737));
  NOR2_X1   g537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  NOR2_X1   g540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g541(.A1(new_n649), .A2(new_n259), .ZN(new_n742));
  INV_X1    g542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g543(.A(new_n743), .B1(new_n255), .B2(G45), .ZN(new_n744));
  OAI21_X1  g544(.A(new_n744), .B1(G45), .B2(new_n234), .ZN(new_n745));
  INV_X1    g545(.A(G355), .ZN(new_n746));
  NAND2_X1  g546(.A1(new_n259), .A2(new_n236), .ZN(new_n747));
  OAI221_X1 g547(.A(new_n745), .B1(G116), .B2(new_n236), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI22_X1  g548(.A1(new_n735), .A2(new_n737), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  INV_X1    g549(.A(new_n740), .ZN(new_n750));
  OAI21_X1  g550(.A(new_n749), .B1(new_n640), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g551(.A(new_n688), .B1(new_n689), .B2(new_n751), .ZN(G396));
  NOR2_X1   g552(.A1(new_n428), .A2(new_n630), .ZN(new_n753));
  NAND2_X1  g553(.A1(new_n351), .A2(new_n630), .ZN(new_n754));
  NAND2_X1  g554(.A1(new_n362), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n428), .ZN(new_n756));
  INV_X1    g556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g557(.A1(new_n664), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g558(.A1(new_n601), .A2(new_n616), .A3(new_n618), .ZN(new_n759));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n631), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g561(.A(new_n680), .ZN(new_n762));
  XNOR2_X1  g562(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n689), .ZN(new_n764));
  AOI21_X1  g564(.A(new_n689), .B1(new_n757), .B2(new_n738), .ZN(new_n765));
  NOR2_X1   g565(.A1(new_n737), .A2(new_n738), .ZN(new_n766));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n298), .ZN(new_n767));
  AOI22_X1  g567(.A1(new_n704), .A2(G116), .B1(G303), .B2(new_n697), .ZN(new_n768));
  OR2_X1    g568(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g569(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n770));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g571(.A(G283), .ZN(new_n772));
  OAI21_X1  g572(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g573(.A(new_n773), .B(KEYINPUT98), .ZN(new_n774));
  OAI211_X1 g574(.A(new_n774), .B(new_n325), .C1(new_n219), .C2(new_n714), .ZN(new_n775));
  OAI22_X1  g575(.A1(new_n694), .A2(new_n702), .B1(new_n211), .B2(new_n719), .ZN(new_n776));
  INV_X1    g576(.A(new_n701), .ZN(new_n777));
  AOI22_X1  g577(.A1(new_n717), .A2(G294), .B1(new_n777), .B2(G97), .ZN(new_n778));
  XOR2_X1   g578(.A(new_n778), .B(KEYINPUT99), .Z(new_n779));
  NOR3_X1   g579(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g580(.A1(new_n720), .A2(G68), .ZN(new_n781));
  INV_X1    g581(.A(G132), .ZN(new_n782));
  AOI22_X1  g582(.A1(new_n707), .A2(G150), .B1(G143), .B2(new_n717), .ZN(new_n783));
  INV_X1    g583(.A(G137), .ZN(new_n784));
  OAI221_X1 g584(.A(new_n783), .B1(new_n784), .B2(new_n723), .C1(new_n728), .C2(new_n705), .ZN(new_n785));
  INV_X1    g585(.A(KEYINPUT34), .ZN(new_n786));
  OAI221_X1 g586(.A(new_n781), .B1(new_n782), .B2(new_n694), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g587(.A(new_n325), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g588(.A(new_n788), .B1(new_n202), .B2(new_n714), .ZN(new_n789));
  AOI211_X1 g589(.A(new_n787), .B(new_n789), .C1(G58), .C2(new_n777), .ZN(new_n790));
  OAI21_X1  g590(.A(new_n737), .B1(new_n780), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g591(.A1(new_n765), .A2(new_n767), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g592(.A1(new_n764), .A2(new_n792), .ZN(G384));
  NOR2_X1   g593(.A1(new_n315), .A2(new_n630), .ZN(new_n794));
  INV_X1    g594(.A(new_n628), .ZN(new_n795));
  NAND2_X1  g595(.A1(new_n400), .A2(new_n795), .ZN(new_n796));
  INV_X1    g596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g597(.A(new_n797), .B1(new_n418), .B2(new_n425), .ZN(new_n798));
  AND3_X1   g598(.A1(new_n379), .A2(new_n398), .A3(new_n392), .ZN(new_n799));
  AOI21_X1  g599(.A(new_n398), .B1(new_n379), .B2(new_n392), .ZN(new_n800));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n800), .A3(new_n396), .ZN(new_n801));
  OAI21_X1  g601(.A(new_n423), .B1(new_n801), .B2(new_n628), .ZN(new_n802));
  NOR2_X1   g602(.A1(new_n801), .A2(new_n414), .ZN(new_n803));
  OAI21_X1  g603(.A(KEYINPUT37), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g604(.A1(new_n400), .A2(new_n415), .ZN(new_n805));
  INV_X1    g605(.A(KEYINPUT37), .ZN(new_n806));
  NAND4_X1  g606(.A1(new_n805), .A2(new_n796), .A3(new_n806), .A4(new_n423), .ZN(new_n807));
  NAND3_X1  g607(.A1(new_n804), .A2(KEYINPUT104), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g608(.A1(new_n802), .A2(new_n803), .ZN(new_n809));
  INV_X1    g609(.A(KEYINPUT104), .ZN(new_n810));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n806), .ZN(new_n811));
  NAND3_X1  g611(.A1(new_n798), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  INV_X1    g612(.A(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n815));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g616(.A(KEYINPUT39), .ZN(new_n817));
  OAI21_X1  g617(.A(new_n365), .B1(new_n377), .B2(new_n378), .ZN(new_n818));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n391), .ZN(new_n819));
  INV_X1    g619(.A(KEYINPUT103), .ZN(new_n820));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n820), .A3(new_n302), .ZN(new_n821));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n379), .ZN(new_n822));
  AOI21_X1  g622(.A(new_n820), .B1(new_n819), .B2(new_n302), .ZN(new_n823));
  OAI21_X1  g623(.A(new_n397), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g624(.A(new_n795), .B(new_n824), .C1(new_n418), .C2(new_n425), .ZN(new_n825));
  NAND2_X1  g625(.A1(new_n414), .A2(new_n628), .ZN(new_n826));
  AOI22_X1  g626(.A1(new_n824), .A2(new_n826), .B1(new_n422), .B2(new_n801), .ZN(new_n827));
  OAI21_X1  g627(.A(new_n807), .B1(new_n827), .B2(new_n806), .ZN(new_n828));
  NAND3_X1  g628(.A1(new_n825), .A2(KEYINPUT38), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g629(.A1(new_n812), .A2(KEYINPUT105), .A3(new_n813), .ZN(new_n830));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n817), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g631(.A(KEYINPUT106), .ZN(new_n832));
  INV_X1    g632(.A(new_n829), .ZN(new_n833));
  AOI21_X1  g633(.A(KEYINPUT38), .B1(new_n825), .B2(new_n828), .ZN(new_n834));
  OAI21_X1  g634(.A(KEYINPUT39), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g635(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g636(.A(new_n832), .B1(new_n831), .B2(new_n835), .ZN(new_n837));
  OAI21_X1  g637(.A(new_n794), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g638(.A1(new_n593), .A2(new_n795), .ZN(new_n839));
  INV_X1    g639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g640(.A1(new_n314), .A2(new_n630), .ZN(new_n841));
  NAND3_X1  g641(.A1(new_n315), .A2(new_n343), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g642(.A1(new_n294), .A2(new_n314), .A3(new_n630), .ZN(new_n843));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g644(.A(new_n844), .ZN(new_n845));
  INV_X1    g645(.A(new_n753), .ZN(new_n846));
  AOI21_X1  g646(.A(new_n845), .B1(new_n760), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g647(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  OAI21_X1  g648(.A(new_n848), .B1(new_n834), .B2(new_n833), .ZN(new_n849));
  NAND3_X1  g649(.A1(new_n838), .A2(new_n840), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g650(.A(new_n850), .B(KEYINPUT108), .Z(new_n851));
  OAI21_X1  g651(.A(new_n429), .B1(new_n663), .B2(new_n665), .ZN(new_n852));
  AND2_X1   g652(.A1(new_n852), .A2(new_n597), .ZN(new_n853));
  XNOR2_X1  g653(.A(new_n851), .B(new_n853), .ZN(new_n854));
  NAND4_X1  g654(.A1(new_n677), .A2(new_n844), .A3(new_n678), .A4(new_n756), .ZN(new_n855));
  INV_X1    g655(.A(new_n834), .ZN(new_n856));
  AOI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n829), .ZN(new_n857));
  OAI21_X1  g657(.A(KEYINPUT107), .B1(new_n857), .B2(KEYINPUT40), .ZN(new_n858));
  INV_X1    g658(.A(KEYINPUT107), .ZN(new_n859));
  INV_X1    g659(.A(KEYINPUT40), .ZN(new_n860));
  NOR2_X1   g660(.A1(new_n833), .A2(new_n834), .ZN(new_n861));
  OAI211_X1 g661(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n855), .ZN(new_n862));
  NAND2_X1  g662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g663(.A1(new_n816), .A2(new_n829), .A3(new_n830), .ZN(new_n864));
  INV_X1    g664(.A(new_n855), .ZN(new_n865));
  NAND3_X1  g665(.A1(new_n864), .A2(KEYINPUT40), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g666(.A1(new_n863), .A2(new_n429), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g667(.A1(new_n863), .A2(G330), .A3(new_n866), .ZN(new_n868));
  NAND2_X1  g668(.A1(new_n762), .A2(new_n429), .ZN(new_n869));
  AOI22_X1  g669(.A1(new_n867), .A2(new_n679), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g670(.A(new_n854), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g671(.A(new_n871), .B1(new_n272), .B2(new_n624), .ZN(new_n872));
  OAI21_X1  g672(.A(G77), .B1(new_n217), .B2(new_n222), .ZN(new_n873));
  OAI22_X1  g673(.A1(new_n873), .A2(new_n234), .B1(G50), .B2(new_n222), .ZN(new_n874));
  NAND3_X1  g674(.A1(new_n874), .A2(G1), .A3(new_n623), .ZN(new_n875));
  XOR2_X1   g675(.A(new_n875), .B(KEYINPUT101), .Z(new_n876));
  INV_X1    g676(.A(KEYINPUT35), .ZN(new_n877));
  AOI211_X1 g677(.A(new_n233), .B(new_n232), .C1(new_n535), .C2(new_n877), .ZN(new_n878));
  OAI211_X1 g678(.A(new_n878), .B(G116), .C1(new_n877), .C2(new_n535), .ZN(new_n879));
  XOR2_X1   g679(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n880));
  XNOR2_X1  g680(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND3_X1  g681(.A1(new_n872), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  XOR2_X1   g682(.A(new_n882), .B(KEYINPUT109), .Z(G367));
  OAI21_X1  g683(.A(new_n644), .B1(new_n641), .B2(new_n635), .ZN(new_n884));
  NOR2_X1   g684(.A1(new_n681), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g685(.A1(new_n643), .A2(new_n646), .ZN(new_n886));
  OAI211_X1 g686(.A(new_n551), .B(new_n554), .C1(new_n539), .C2(new_n631), .ZN(new_n887));
  OAI21_X1  g687(.A(new_n887), .B1(new_n554), .B2(new_n631), .ZN(new_n888));
  INV_X1    g688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g690(.A(new_n890), .B(KEYINPUT44), .Z(new_n891));
  NOR2_X1   g691(.A1(new_n886), .A2(new_n889), .ZN(new_n892));
  XNOR2_X1  g692(.A(new_n892), .B(KEYINPUT45), .ZN(new_n893));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g694(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n682), .ZN(new_n896));
  XNOR2_X1  g696(.A(new_n650), .B(KEYINPUT41), .ZN(new_n897));
  AOI21_X1  g697(.A(new_n686), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g698(.A1(new_n643), .A2(new_n887), .ZN(new_n899));
  XNOR2_X1  g699(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  OAI21_X1  g700(.A(new_n554), .B1(new_n887), .B2(new_n589), .ZN(new_n901));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n631), .ZN(new_n902));
  OR2_X1    g702(.A1(new_n631), .A2(new_n562), .ZN(new_n903));
  NAND2_X1  g703(.A1(new_n584), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g704(.A(new_n904), .B1(new_n583), .B2(new_n903), .ZN(new_n905));
  AOI22_X1  g705(.A1(new_n900), .A2(new_n902), .B1(KEYINPUT43), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g706(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n907));
  XNOR2_X1  g707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NOR2_X1   g708(.A1(new_n642), .A2(new_n889), .ZN(new_n909));
  XNOR2_X1  g709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g710(.A1(new_n905), .A2(new_n750), .ZN(new_n911));
  OAI221_X1 g711(.A(new_n741), .B1(new_n236), .B2(new_n348), .C1(new_n247), .C2(new_n743), .ZN(new_n912));
  XNOR2_X1  g712(.A(new_n912), .B(KEYINPUT111), .ZN(new_n913));
  AOI22_X1  g713(.A1(new_n704), .A2(G283), .B1(G311), .B2(new_n697), .ZN(new_n914));
  NAND2_X1  g714(.A1(new_n720), .A2(G97), .ZN(new_n915));
  NAND2_X1  g715(.A1(new_n777), .A2(G107), .ZN(new_n916));
  AOI21_X1  g716(.A(new_n259), .B1(new_n717), .B2(G303), .ZN(new_n917));
  NAND4_X1  g717(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g718(.A1(new_n695), .A2(G317), .ZN(new_n919));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n920));
  NAND2_X1  g720(.A1(new_n715), .A2(G116), .ZN(new_n921));
  OAI221_X1 g721(.A(new_n919), .B1(new_n920), .B2(new_n921), .C1(new_n699), .C2(new_n771), .ZN(new_n922));
  AOI211_X1 g722(.A(new_n918), .B(new_n922), .C1(new_n920), .C2(new_n921), .ZN(new_n923));
  NAND2_X1  g723(.A1(new_n704), .A2(G50), .ZN(new_n924));
  INV_X1    g724(.A(new_n771), .ZN(new_n925));
  AOI22_X1  g725(.A1(new_n925), .A2(G159), .B1(G150), .B2(new_n717), .ZN(new_n926));
  OAI21_X1  g726(.A(new_n926), .B1(new_n222), .B2(new_n701), .ZN(new_n927));
  OAI21_X1  g727(.A(new_n259), .B1(new_n694), .B2(new_n784), .ZN(new_n928));
  NAND2_X1  g728(.A1(new_n697), .A2(G143), .ZN(new_n929));
  OAI221_X1 g729(.A(new_n929), .B1(new_n298), .B2(new_n719), .C1(new_n714), .C2(new_n217), .ZN(new_n930));
  NOR3_X1   g730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g731(.A(new_n923), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g732(.A(new_n932), .B(KEYINPUT47), .ZN(new_n933));
  INV_X1    g733(.A(new_n737), .ZN(new_n934));
  OAI211_X1 g734(.A(new_n687), .B(new_n913), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OAI22_X1  g735(.A1(new_n898), .A2(new_n910), .B1(new_n911), .B2(new_n935), .ZN(G387));
  OAI21_X1  g736(.A(new_n742), .B1(new_n244), .B2(new_n280), .ZN(new_n937));
  OAI21_X1  g737(.A(new_n937), .B1(new_n653), .B2(new_n747), .ZN(new_n938));
  OAI211_X1 g738(.A(new_n653), .B(new_n280), .C1(new_n222), .C2(new_n298), .ZN(new_n939));
  NAND2_X1  g739(.A1(new_n319), .A2(new_n202), .ZN(new_n940));
  XNOR2_X1  g740(.A(new_n940), .B(KEYINPUT50), .ZN(new_n941));
  OAI21_X1  g741(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g742(.A1(new_n649), .A2(new_n219), .ZN(new_n943));
  AOI211_X1 g743(.A(new_n740), .B(new_n737), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  OAI221_X1 g744(.A(new_n259), .B1(new_n222), .B2(new_n705), .C1(new_n694), .C2(new_n317), .ZN(new_n945));
  AOI21_X1  g745(.A(new_n945), .B1(new_n319), .B2(new_n707), .ZN(new_n946));
  NOR2_X1   g746(.A1(new_n701), .A2(new_n348), .ZN(new_n947));
  NOR2_X1   g747(.A1(new_n714), .A2(new_n298), .ZN(new_n948));
  AOI211_X1 g748(.A(new_n947), .B(new_n948), .C1(G159), .C2(new_n697), .ZN(new_n949));
  NAND2_X1  g749(.A1(new_n717), .A2(G50), .ZN(new_n950));
  NAND4_X1  g750(.A1(new_n946), .A2(new_n915), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  AOI22_X1  g751(.A1(new_n704), .A2(G303), .B1(G317), .B2(new_n717), .ZN(new_n952));
  INV_X1    g752(.A(G322), .ZN(new_n953));
  OAI221_X1 g753(.A(new_n952), .B1(new_n953), .B2(new_n723), .C1(new_n771), .C2(new_n702), .ZN(new_n954));
  XNOR2_X1  g754(.A(new_n954), .B(KEYINPUT48), .ZN(new_n955));
  OAI221_X1 g755(.A(new_n955), .B1(new_n772), .B2(new_n701), .C1(new_n699), .C2(new_n714), .ZN(new_n956));
  XOR2_X1   g756(.A(new_n956), .B(KEYINPUT49), .Z(new_n957));
  NAND2_X1  g757(.A1(new_n695), .A2(G326), .ZN(new_n958));
  AOI21_X1  g758(.A(new_n259), .B1(new_n720), .B2(G116), .ZN(new_n959));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g760(.A(new_n951), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  AOI211_X1 g761(.A(new_n689), .B(new_n944), .C1(new_n961), .C2(new_n737), .ZN(new_n962));
  OAI21_X1  g762(.A(new_n962), .B1(new_n633), .B2(new_n750), .ZN(new_n963));
  INV_X1    g763(.A(new_n884), .ZN(new_n964));
  OAI21_X1  g764(.A(new_n650), .B1(new_n682), .B2(new_n964), .ZN(new_n965));
  OAI221_X1 g765(.A(new_n963), .B1(new_n685), .B2(new_n884), .C1(new_n965), .C2(new_n885), .ZN(G393));
  XOR2_X1   g766(.A(new_n894), .B(new_n642), .Z(new_n967));
  OAI21_X1  g767(.A(new_n967), .B1(new_n681), .B2(new_n884), .ZN(new_n968));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n650), .A3(new_n895), .ZN(new_n969));
  AOI22_X1  g769(.A1(new_n925), .A2(G303), .B1(G116), .B2(new_n777), .ZN(new_n970));
  NAND2_X1  g770(.A1(new_n695), .A2(G322), .ZN(new_n971));
  OAI21_X1  g771(.A(new_n732), .B1(new_n772), .B2(new_n714), .ZN(new_n972));
  AOI211_X1 g772(.A(new_n259), .B(new_n972), .C1(G294), .C2(new_n704), .ZN(new_n973));
  AOI22_X1  g773(.A1(G311), .A2(new_n717), .B1(new_n697), .B2(G317), .ZN(new_n974));
  XOR2_X1   g774(.A(new_n974), .B(KEYINPUT52), .Z(new_n975));
  NAND4_X1  g775(.A1(new_n970), .A2(new_n971), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g776(.A1(new_n771), .A2(new_n202), .B1(new_n320), .B2(new_n705), .ZN(new_n977));
  XOR2_X1   g777(.A(new_n977), .B(KEYINPUT113), .Z(new_n978));
  OAI221_X1 g778(.A(new_n259), .B1(new_n211), .B2(new_n719), .C1(new_n714), .C2(new_n222), .ZN(new_n979));
  AOI21_X1  g779(.A(new_n979), .B1(new_n695), .B2(G143), .ZN(new_n980));
  XOR2_X1   g780(.A(new_n980), .B(KEYINPUT112), .Z(new_n981));
  INV_X1    g781(.A(new_n717), .ZN(new_n982));
  OAI22_X1  g782(.A1(new_n317), .A2(new_n723), .B1(new_n982), .B2(new_n728), .ZN(new_n983));
  INV_X1    g783(.A(KEYINPUT51), .ZN(new_n984));
  AOI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(G77), .B2(new_n777), .ZN(new_n985));
  NAND3_X1  g785(.A1(new_n978), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g786(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  OAI21_X1  g787(.A(new_n976), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n737), .ZN(new_n989));
  NAND2_X1  g789(.A1(new_n889), .A2(new_n740), .ZN(new_n990));
  OAI221_X1 g790(.A(new_n741), .B1(new_n436), .B2(new_n236), .C1(new_n252), .C2(new_n743), .ZN(new_n991));
  NAND4_X1  g791(.A1(new_n989), .A2(new_n990), .A3(new_n687), .A4(new_n991), .ZN(new_n992));
  OAI211_X1 g792(.A(new_n969), .B(new_n992), .C1(new_n685), .C2(new_n967), .ZN(G390));
  NAND4_X1  g793(.A1(new_n677), .A2(new_n678), .A3(G330), .A4(new_n756), .ZN(new_n994));
  OR2_X1    g794(.A1(new_n994), .A2(new_n845), .ZN(new_n995));
  INV_X1    g795(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g796(.A1(new_n760), .A2(new_n846), .ZN(new_n997));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n844), .ZN(new_n998));
  INV_X1    g798(.A(KEYINPUT114), .ZN(new_n999));
  INV_X1    g799(.A(new_n794), .ZN(new_n1000));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g801(.A(KEYINPUT114), .B1(new_n847), .B2(new_n794), .ZN(new_n1002));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g803(.A1(new_n836), .A2(new_n1003), .A3(new_n837), .ZN(new_n1004));
  INV_X1    g804(.A(new_n864), .ZN(new_n1005));
  AOI21_X1  g805(.A(new_n753), .B1(new_n662), .B2(new_n362), .ZN(new_n1006));
  OAI21_X1  g806(.A(new_n1000), .B1(new_n1006), .B2(new_n845), .ZN(new_n1007));
  NOR2_X1   g807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g808(.A(new_n996), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g809(.A(new_n1008), .ZN(new_n1010));
  INV_X1    g810(.A(new_n837), .ZN(new_n1011));
  NAND3_X1  g811(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n1012));
  NAND2_X1  g812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g813(.A(new_n995), .B(new_n1010), .C1(new_n1013), .C2(new_n1003), .ZN(new_n1014));
  NAND3_X1  g814(.A1(new_n1009), .A2(new_n1014), .A3(new_n686), .ZN(new_n1015));
  NAND2_X1  g815(.A1(new_n766), .A2(new_n320), .ZN(new_n1016));
  NOR2_X1   g816(.A1(new_n714), .A2(new_n317), .ZN(new_n1017));
  XNOR2_X1  g817(.A(new_n1017), .B(KEYINPUT53), .ZN(new_n1018));
  INV_X1    g818(.A(G128), .ZN(new_n1019));
  OAI221_X1 g819(.A(new_n1018), .B1(new_n1019), .B2(new_n723), .C1(new_n728), .C2(new_n701), .ZN(new_n1020));
  AOI22_X1  g820(.A1(new_n925), .A2(G137), .B1(G125), .B2(new_n695), .ZN(new_n1021));
  XOR2_X1   g821(.A(KEYINPUT54), .B(G143), .Z(new_n1022));
  XNOR2_X1  g822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  AOI21_X1  g823(.A(new_n325), .B1(new_n704), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g824(.A(new_n1021), .B(new_n1024), .C1(new_n782), .C2(new_n982), .ZN(new_n1025));
  AOI211_X1 g825(.A(new_n1020), .B(new_n1025), .C1(G50), .C2(new_n720), .ZN(new_n1026));
  XNOR2_X1  g826(.A(new_n1026), .B(KEYINPUT117), .ZN(new_n1027));
  OAI221_X1 g827(.A(new_n781), .B1(new_n772), .B2(new_n723), .C1(new_n694), .C2(new_n699), .ZN(new_n1028));
  OAI22_X1  g828(.A1(new_n714), .A2(new_n211), .B1(new_n298), .B2(new_n701), .ZN(new_n1029));
  NOR2_X1   g829(.A1(new_n982), .A2(new_n213), .ZN(new_n1030));
  NOR4_X1   g830(.A1(new_n1028), .A2(new_n259), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI221_X1 g831(.A(new_n1031), .B1(new_n436), .B2(new_n705), .C1(new_n219), .C2(new_n771), .ZN(new_n1032));
  NAND2_X1  g832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g833(.A(new_n1033), .B(KEYINPUT118), .ZN(new_n1034));
  AOI21_X1  g834(.A(new_n689), .B1(new_n1034), .B2(new_n737), .ZN(new_n1035));
  OAI211_X1 g835(.A(new_n1016), .B(new_n1035), .C1(new_n1013), .C2(new_n739), .ZN(new_n1036));
  NAND2_X1  g836(.A1(new_n1015), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g837(.A1(new_n994), .A2(new_n845), .ZN(new_n1038));
  NAND2_X1  g838(.A1(new_n995), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g839(.A1(new_n1039), .A2(new_n997), .ZN(new_n1040));
  NAND3_X1  g840(.A1(new_n995), .A2(new_n1006), .A3(new_n1038), .ZN(new_n1041));
  NAND2_X1  g841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AND4_X1   g842(.A1(new_n597), .A2(new_n1042), .A3(new_n852), .A4(new_n869), .ZN(new_n1043));
  AOI21_X1  g843(.A(new_n1043), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1044));
  NAND3_X1  g844(.A1(new_n1009), .A2(new_n1014), .A3(new_n1043), .ZN(new_n1045));
  INV_X1    g845(.A(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g847(.A1(new_n1009), .A2(new_n1014), .A3(KEYINPUT115), .A4(new_n1043), .ZN(new_n1048));
  AOI21_X1  g848(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g849(.A(new_n1037), .B1(new_n1049), .B2(new_n650), .ZN(new_n1050));
  INV_X1    g850(.A(new_n1050), .ZN(G378));
  OAI22_X1  g851(.A1(new_n705), .A2(new_n348), .B1(new_n222), .B2(new_n701), .ZN(new_n1052));
  NOR3_X1   g852(.A1(new_n948), .A2(new_n648), .A3(new_n259), .ZN(new_n1053));
  XNOR2_X1  g853(.A(new_n1053), .B(KEYINPUT119), .ZN(new_n1054));
  OAI221_X1 g854(.A(new_n1054), .B1(new_n217), .B2(new_n719), .C1(new_n772), .C2(new_n694), .ZN(new_n1055));
  XOR2_X1   g855(.A(new_n1055), .B(KEYINPUT120), .Z(new_n1056));
  AOI211_X1 g856(.A(new_n1052), .B(new_n1056), .C1(G107), .C2(new_n717), .ZN(new_n1057));
  OAI221_X1 g857(.A(new_n1057), .B1(new_n436), .B2(new_n725), .C1(new_n213), .C2(new_n723), .ZN(new_n1058));
  XNOR2_X1  g858(.A(new_n1058), .B(KEYINPUT58), .ZN(new_n1059));
  AOI22_X1  g859(.A1(G132), .A2(new_n707), .B1(new_n704), .B2(G137), .ZN(new_n1060));
  AOI22_X1  g860(.A1(new_n715), .A2(new_n1023), .B1(new_n717), .B2(G128), .ZN(new_n1061));
  NAND2_X1  g861(.A1(new_n777), .A2(G150), .ZN(new_n1062));
  NAND2_X1  g862(.A1(new_n697), .A2(G125), .ZN(new_n1063));
  NAND4_X1  g863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  XOR2_X1   g864(.A(new_n1064), .B(KEYINPUT59), .Z(new_n1065));
  AOI211_X1 g865(.A(G33), .B(G41), .C1(new_n695), .C2(G124), .ZN(new_n1066));
  OAI211_X1 g866(.A(new_n1065), .B(new_n1066), .C1(new_n728), .C2(new_n719), .ZN(new_n1067));
  OAI221_X1 g867(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n648), .C2(new_n259), .ZN(new_n1068));
  NAND3_X1  g868(.A1(new_n1059), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g869(.A(new_n1069), .B(KEYINPUT121), .ZN(new_n1070));
  NAND2_X1  g870(.A1(new_n1070), .A2(new_n737), .ZN(new_n1071));
  NAND2_X1  g871(.A1(new_n323), .A2(new_n795), .ZN(new_n1072));
  XNOR2_X1  g872(.A(new_n340), .B(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g873(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1074));
  XNOR2_X1  g874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  NAND2_X1  g875(.A1(new_n1075), .A2(new_n738), .ZN(new_n1076));
  NAND2_X1  g876(.A1(new_n766), .A2(new_n202), .ZN(new_n1077));
  NAND4_X1  g877(.A1(new_n1071), .A2(new_n687), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g878(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g879(.A(KEYINPUT122), .ZN(new_n1080));
  NAND4_X1  g880(.A1(new_n863), .A2(new_n1080), .A3(G330), .A4(new_n866), .ZN(new_n1081));
  INV_X1    g881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g882(.A1(new_n850), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g883(.A1(new_n1081), .A2(new_n838), .A3(new_n840), .A4(new_n849), .ZN(new_n1084));
  AOI21_X1  g884(.A(new_n1075), .B1(new_n868), .B2(KEYINPUT122), .ZN(new_n1085));
  AND3_X1   g885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g886(.A(new_n1085), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1087));
  NOR2_X1   g887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g888(.A(new_n1079), .B1(new_n1088), .B2(new_n686), .ZN(new_n1089));
  NAND2_X1  g889(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1090));
  NAND2_X1  g890(.A1(new_n853), .A2(new_n869), .ZN(new_n1091));
  INV_X1    g891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g893(.A(KEYINPUT57), .B1(new_n1093), .B2(new_n1088), .ZN(new_n1094));
  AOI21_X1  g894(.A(new_n1091), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1095));
  NAND2_X1  g895(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1096));
  INV_X1    g896(.A(new_n1085), .ZN(new_n1097));
  NAND2_X1  g897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g898(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1099));
  NAND3_X1  g899(.A1(new_n1098), .A2(KEYINPUT57), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g900(.A(new_n650), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g901(.A(new_n1089), .B1(new_n1094), .B2(new_n1101), .ZN(G375));
  INV_X1    g902(.A(new_n1042), .ZN(new_n1103));
  NAND2_X1  g903(.A1(new_n1091), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g904(.A(new_n1043), .ZN(new_n1105));
  NAND3_X1  g905(.A1(new_n1104), .A2(new_n897), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g906(.A(new_n689), .B1(new_n845), .B2(new_n738), .ZN(new_n1107));
  OAI221_X1 g907(.A(new_n259), .B1(new_n782), .B2(new_n723), .C1(new_n705), .C2(new_n317), .ZN(new_n1108));
  OAI22_X1  g908(.A1(new_n694), .A2(new_n1019), .B1(new_n728), .B2(new_n714), .ZN(new_n1109));
  XOR2_X1   g909(.A(new_n1109), .B(KEYINPUT123), .Z(new_n1110));
  AOI22_X1  g910(.A1(new_n720), .A2(G58), .B1(G50), .B2(new_n777), .ZN(new_n1111));
  OAI211_X1 g911(.A(new_n1110), .B(new_n1111), .C1(new_n784), .C2(new_n982), .ZN(new_n1112));
  AOI211_X1 g912(.A(new_n1108), .B(new_n1112), .C1(new_n925), .C2(new_n1023), .ZN(new_n1113));
  AOI22_X1  g913(.A1(new_n925), .A2(G116), .B1(G294), .B2(new_n697), .ZN(new_n1114));
  OAI221_X1 g914(.A(new_n1114), .B1(new_n436), .B2(new_n714), .C1(new_n219), .C2(new_n705), .ZN(new_n1115));
  AND2_X1   g915(.A1(new_n695), .A2(G303), .ZN(new_n1116));
  OAI221_X1 g916(.A(new_n325), .B1(new_n298), .B2(new_n719), .C1(new_n982), .C2(new_n772), .ZN(new_n1117));
  NOR4_X1   g917(.A1(new_n1115), .A2(new_n947), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g918(.A(new_n737), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g919(.A1(new_n1107), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g920(.A(new_n1120), .B1(new_n222), .B2(new_n766), .ZN(new_n1121));
  AOI21_X1  g921(.A(new_n1121), .B1(new_n1042), .B2(new_n686), .ZN(new_n1122));
  NAND2_X1  g922(.A1(new_n1106), .A2(new_n1122), .ZN(G381));
  INV_X1    g923(.A(KEYINPUT57), .ZN(new_n1124));
  NOR3_X1   g924(.A1(new_n1086), .A2(new_n1087), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g925(.A1(new_n1093), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g926(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1127));
  OAI21_X1  g927(.A(new_n1124), .B1(new_n1095), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g928(.A1(new_n1126), .A2(new_n1128), .A3(new_n650), .ZN(new_n1129));
  NAND3_X1  g929(.A1(new_n1129), .A2(new_n1050), .A3(new_n1089), .ZN(new_n1130));
  NOR3_X1   g930(.A1(new_n1130), .A2(G384), .A3(G381), .ZN(new_n1131));
  OR2_X1    g931(.A1(G387), .A2(G390), .ZN(new_n1132));
  NOR3_X1   g932(.A1(new_n1132), .A2(G396), .A3(G393), .ZN(new_n1133));
  NAND2_X1  g933(.A1(new_n1131), .A2(new_n1133), .ZN(G407));
  OAI211_X1 g934(.A(G407), .B(G213), .C1(G343), .C2(new_n1130), .ZN(G409));
  OAI21_X1  g935(.A(KEYINPUT124), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1136));
  INV_X1    g936(.A(KEYINPUT124), .ZN(new_n1137));
  NAND3_X1  g937(.A1(new_n1098), .A2(new_n1137), .A3(new_n1099), .ZN(new_n1138));
  NAND3_X1  g938(.A1(new_n1136), .A2(new_n1138), .A3(new_n686), .ZN(new_n1139));
  AND2_X1   g939(.A1(new_n1050), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g940(.A1(new_n1095), .A2(new_n1127), .ZN(new_n1141));
  AOI21_X1  g941(.A(new_n1079), .B1(new_n1141), .B2(new_n897), .ZN(new_n1142));
  AOI22_X1  g942(.A1(new_n1140), .A2(new_n1142), .B1(G213), .B2(new_n629), .ZN(new_n1143));
  NAND2_X1  g943(.A1(G375), .A2(G378), .ZN(new_n1144));
  NAND2_X1  g944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g945(.A(KEYINPUT60), .ZN(new_n1146));
  AOI21_X1  g946(.A(new_n651), .B1(new_n1104), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g947(.A(new_n1147), .B(new_n1105), .C1(new_n1146), .C2(new_n1104), .ZN(new_n1148));
  NAND2_X1  g948(.A1(new_n1148), .A2(new_n1122), .ZN(new_n1149));
  INV_X1    g949(.A(G384), .ZN(new_n1150));
  NAND2_X1  g950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g951(.A1(new_n1148), .A2(new_n1122), .A3(G384), .ZN(new_n1152));
  NAND2_X1  g952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g953(.A1(new_n629), .A2(G213), .A3(G2897), .ZN(new_n1154));
  XNOR2_X1  g954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AOI21_X1  g955(.A(KEYINPUT61), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g956(.A(new_n1050), .B1(new_n1129), .B2(new_n1089), .ZN(new_n1157));
  NAND3_X1  g957(.A1(new_n1093), .A2(new_n897), .A3(new_n1088), .ZN(new_n1158));
  NAND4_X1  g958(.A1(new_n1158), .A2(new_n1050), .A3(new_n1078), .A4(new_n1139), .ZN(new_n1159));
  NAND2_X1  g959(.A1(new_n629), .A2(G213), .ZN(new_n1160));
  NAND2_X1  g960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g961(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g962(.A(new_n1153), .ZN(new_n1163));
  AOI21_X1  g963(.A(KEYINPUT62), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND4_X1   g964(.A1(KEYINPUT62), .A2(new_n1143), .A3(new_n1163), .A4(new_n1144), .ZN(new_n1165));
  OAI21_X1  g965(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g966(.A(KEYINPUT127), .ZN(new_n1167));
  NAND2_X1  g967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g968(.A(G393), .B(G396), .ZN(new_n1169));
  NAND2_X1  g969(.A1(G387), .A2(G390), .ZN(new_n1170));
  AND3_X1   g970(.A1(new_n1132), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g971(.A(new_n1169), .B1(new_n1132), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g973(.A(new_n1173), .ZN(new_n1174));
  OAI211_X1 g974(.A(new_n1156), .B(KEYINPUT127), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1175));
  NAND3_X1  g975(.A1(new_n1168), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g976(.A(KEYINPUT63), .ZN(new_n1177));
  OAI21_X1  g977(.A(new_n1177), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1178));
  INV_X1    g978(.A(KEYINPUT125), .ZN(new_n1179));
  NAND2_X1  g979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g980(.A(KEYINPUT125), .B(new_n1177), .C1(new_n1145), .C2(new_n1153), .ZN(new_n1181));
  NAND2_X1  g981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g982(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1183));
  AOI21_X1  g983(.A(KEYINPUT61), .B1(new_n1183), .B2(KEYINPUT63), .ZN(new_n1184));
  OR2_X1    g984(.A1(new_n1145), .A2(KEYINPUT126), .ZN(new_n1185));
  NAND2_X1  g985(.A1(new_n1145), .A2(KEYINPUT126), .ZN(new_n1186));
  NAND3_X1  g986(.A1(new_n1185), .A2(new_n1155), .A3(new_n1186), .ZN(new_n1187));
  NAND4_X1  g987(.A1(new_n1182), .A2(new_n1184), .A3(new_n1173), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g988(.A1(new_n1176), .A2(new_n1188), .ZN(G405));
  NAND2_X1  g989(.A1(new_n1144), .A2(new_n1130), .ZN(new_n1190));
  XNOR2_X1  g990(.A(new_n1190), .B(new_n1163), .ZN(new_n1191));
  XNOR2_X1  g991(.A(new_n1191), .B(new_n1173), .ZN(G402));
endmodule


