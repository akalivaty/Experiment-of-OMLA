//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1209, new_n1210, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n214), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n217), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n212), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n206), .A2(new_n207), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n211), .A2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n230), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n253), .B2(KEYINPUT79), .ZN(new_n260));
  INV_X1    g0060(.A(new_n258), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n250), .B(KEYINPUT68), .Z(new_n262));
  AOI22_X1  g0062(.A1(new_n254), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G87), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G226), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n264), .B1(new_n266), .B2(new_n267), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n230), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(new_n272), .B2(new_n230), .ZN(new_n276));
  INV_X1    g0076(.A(new_n230), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G232), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(G274), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n281), .B(KEYINPUT66), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n274), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n274), .A2(new_n284), .A3(new_n287), .A4(G190), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT76), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT7), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n265), .B2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT3), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n299));
  OAI211_X1 g0099(.A(KEYINPUT7), .B(new_n212), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n202), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G58), .A2(G68), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n203), .A2(new_n205), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n212), .A2(new_n298), .A3(KEYINPUT69), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT69), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G20), .B2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G159), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n293), .B1(new_n311), .B2(KEYINPUT16), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT16), .ZN(new_n313));
  NOR4_X1   g0113(.A1(new_n301), .A2(new_n310), .A3(KEYINPUT76), .A4(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n256), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n313), .B1(new_n301), .B2(new_n310), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT77), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT77), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n313), .C1(new_n301), .C2(new_n310), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n296), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n325), .B2(new_n212), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n294), .B(G20), .C1(new_n323), .C2(new_n324), .ZN(new_n327));
  OAI21_X1  g0127(.A(G68), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n303), .A2(G20), .B1(new_n308), .B2(G159), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n311), .A2(new_n293), .A3(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n257), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n317), .A2(new_n319), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n322), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n263), .B(new_n292), .C1(new_n321), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT17), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n263), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT78), .B1(new_n315), .B2(new_n320), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n333), .A2(new_n334), .A3(new_n322), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT17), .B1(new_n342), .B2(new_n292), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n263), .B1(new_n321), .B2(new_n335), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT80), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(KEYINPUT80), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n288), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(G169), .B2(new_n288), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n347), .A2(new_n348), .A3(new_n352), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n340), .A2(new_n341), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT80), .B1(new_n358), .B2(new_n263), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n346), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n359), .A2(new_n360), .A3(new_n351), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n344), .B(new_n357), .C1(new_n361), .C2(new_n353), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n212), .A2(G33), .ZN(new_n363));
  INV_X1    g0163(.A(G77), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(new_n212), .B2(G68), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT73), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n308), .A2(KEYINPUT74), .A3(G50), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT74), .B1(new_n308), .B2(G50), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n256), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT11), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n261), .A2(new_n202), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n261), .A2(new_n256), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G68), .A3(new_n252), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT75), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n283), .A2(G238), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(G97), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n383), .B1(new_n298), .B2(new_n384), .C1(new_n270), .C2(new_n267), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n273), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n381), .A2(new_n287), .A3(new_n382), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n219), .A2(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n391), .A2(KEYINPUT72), .A3(new_n382), .A4(new_n386), .ZN(new_n392));
  INV_X1    g0192(.A(new_n386), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n390), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n389), .B(new_n392), .C1(new_n382), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(G169), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT13), .B1(new_n393), .B2(new_n390), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n398), .A2(new_n387), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n396), .B1(new_n395), .B2(G169), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n380), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n380), .B1(G190), .B2(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n395), .A2(G200), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n208), .A2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(G150), .ZN(new_n409));
  INV_X1    g0209(.A(new_n308), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n408), .B1(new_n409), .B2(new_n410), .C1(new_n262), .C2(new_n363), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n256), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n207), .B1(new_n211), .B2(G20), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n376), .A2(new_n413), .B1(new_n207), .B2(new_n261), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n265), .A2(G222), .A3(new_n269), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n418), .B1(new_n364), .B2(new_n265), .C1(new_n268), .C2(new_n266), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n273), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n287), .B(new_n420), .C1(new_n267), .C2(new_n282), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n421), .ZN(new_n424));
  OR3_X1    g0224(.A1(new_n417), .A2(KEYINPUT10), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT10), .B1(new_n417), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n421), .A2(G179), .ZN(new_n428));
  INV_X1    g0228(.A(G169), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n428), .A2(new_n415), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT15), .B(G87), .Z(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n435), .A2(new_n363), .B1(new_n212), .B2(new_n364), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n410), .A2(new_n250), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n256), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n252), .A2(G77), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n438), .B1(G77), .B2(new_n258), .C1(new_n259), .C2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT70), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n283), .A2(G244), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n287), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n265), .A2(G232), .A3(new_n269), .ZN(new_n445));
  INV_X1    g0245(.A(G107), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n445), .B1(new_n446), .B2(new_n265), .C1(new_n266), .C2(new_n219), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n273), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G200), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n441), .B(new_n450), .C1(new_n423), .C2(new_n449), .ZN(new_n451));
  INV_X1    g0251(.A(new_n448), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n429), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n453), .A2(new_n440), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n444), .A2(new_n349), .A3(new_n448), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n362), .A2(new_n407), .A3(new_n433), .A4(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n258), .A2(G97), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n376), .B1(G1), .B2(new_n298), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT83), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(KEYINPUT6), .B2(new_n384), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(G20), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n308), .A2(G77), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n446), .B1(new_n295), .B2(new_n300), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n463), .B(new_n256), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(G107), .B1(new_n326), .B2(new_n327), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n469), .A3(new_n470), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n463), .B1(new_n476), .B2(new_n256), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n462), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n211), .A2(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(new_n279), .A3(G274), .A4(new_n276), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  INV_X1    g0286(.A(new_n482), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(new_n480), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(new_n276), .A3(new_n279), .A4(G257), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n265), .A2(G244), .A3(new_n269), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n497), .B2(new_n273), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n349), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n478), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n220), .A2(new_n384), .A3(new_n446), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n504), .A2(new_n298), .A3(new_n384), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(G20), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n384), .B2(new_n363), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n265), .A2(new_n212), .A3(G68), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n257), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n434), .A2(new_n258), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n460), .A2(new_n435), .ZN(new_n512));
  OR3_X1    g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n265), .A2(G244), .A3(G1698), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  OAI221_X1 g0315(.A(new_n514), .B1(new_n298), .B2(new_n515), .C1(new_n270), .C2(new_n219), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n273), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n276), .A2(new_n279), .A3(G274), .A4(new_n486), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n276), .A2(new_n279), .A3(G250), .A4(new_n479), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n429), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n513), .B(new_n524), .C1(G179), .C2(new_n523), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(G200), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n460), .A2(new_n220), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n510), .A2(new_n511), .A3(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n528), .C1(new_n423), .C2(new_n523), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n256), .B1(new_n471), .B2(new_n472), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT83), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n473), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n497), .A2(new_n273), .ZN(new_n533));
  INV_X1    g0333(.A(new_n490), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n498), .A2(G190), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(new_n462), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n502), .A2(new_n525), .A3(new_n529), .A4(new_n538), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n298), .A2(new_n515), .A3(G20), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n212), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n446), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n265), .A2(new_n212), .A3(G87), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT24), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n257), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n549), .B2(new_n548), .ZN(new_n551));
  OR3_X1    g0351(.A1(new_n258), .A2(KEYINPUT25), .A3(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT25), .B1(new_n258), .B2(G107), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(new_n460), .C2(new_n446), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT89), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n558));
  INV_X1    g0358(.A(G294), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n558), .B1(new_n298), .B2(new_n559), .C1(new_n270), .C2(new_n221), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n273), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT90), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n280), .A2(new_n562), .A3(G264), .A4(new_n488), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT91), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n488), .A2(new_n276), .A3(new_n279), .A4(G264), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT90), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n564), .B1(new_n563), .B2(new_n566), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n484), .B(new_n561), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G200), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n561), .A2(new_n484), .ZN(new_n573));
  INV_X1    g0373(.A(new_n566), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n565), .A2(KEYINPUT90), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OR3_X1    g0376(.A1(new_n573), .A2(new_n576), .A3(G190), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n557), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n539), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n495), .B(new_n212), .C1(G33), .C2(new_n384), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n515), .A2(G20), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n256), .A2(KEYINPUT88), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT88), .B1(new_n256), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(KEYINPUT20), .B(new_n581), .C1(new_n583), .C2(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n258), .A2(G116), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n461), .B2(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n488), .A2(new_n276), .A3(new_n279), .A4(G270), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT86), .B1(new_n484), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n484), .A2(KEYINPUT86), .A3(new_n594), .ZN(new_n597));
  INV_X1    g0397(.A(G264), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT87), .B1(new_n266), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT87), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n265), .A2(new_n600), .A3(G264), .A4(G1698), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n265), .A2(G257), .A3(new_n269), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n325), .A2(G303), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n596), .A2(new_n597), .B1(new_n273), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n580), .B1(new_n593), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n592), .A3(G179), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n273), .ZN(new_n608));
  INV_X1    g0408(.A(new_n597), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(new_n595), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n592), .A3(KEYINPUT21), .A4(G169), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT91), .B1(new_n574), .B2(new_n575), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n567), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(G179), .A3(new_n484), .A4(new_n561), .ZN(new_n615));
  OAI21_X1  g0415(.A(G169), .B1(new_n573), .B2(new_n576), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n556), .B2(new_n551), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n592), .B1(new_n610), .B2(G200), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n605), .A2(G190), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n612), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n458), .A2(new_n579), .A3(new_n621), .ZN(G372));
  NOR2_X1   g0422(.A1(new_n342), .A2(new_n351), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT18), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n401), .A2(new_n402), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT92), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n456), .B(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n627), .A2(new_n380), .B1(new_n629), .B2(new_n406), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT93), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n344), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n406), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n633), .A2(new_n631), .A3(new_n403), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n626), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n431), .B1(new_n635), .B2(new_n427), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n579), .B1(new_n617), .B2(new_n612), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n525), .A2(new_n529), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n502), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n638), .B(new_n525), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n637), .B1(new_n458), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n644), .B(KEYINPUT94), .Z(G369));
  NAND3_X1  g0445(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n592), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n612), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n620), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n615), .A2(new_n616), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n557), .ZN(new_n657));
  INV_X1    g0457(.A(new_n651), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n551), .B2(new_n556), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n578), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n617), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n612), .A2(new_n658), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n660), .A3(new_n661), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n661), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT95), .ZN(G399));
  INV_X1    g0469(.A(new_n215), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n211), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n503), .A2(G116), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT96), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n672), .A2(new_n674), .B1(new_n232), .B2(new_n671), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT28), .Z(new_n676));
  NAND2_X1  g0476(.A1(new_n643), .A2(new_n658), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT29), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n658), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n498), .A2(G179), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n570), .A2(new_n681), .A3(new_n523), .A4(new_n610), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n523), .A2(new_n535), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n613), .A2(new_n567), .B1(new_n273), .B2(new_n560), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G179), .A4(new_n605), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n561), .B1(new_n568), .B2(new_n569), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n498), .B(new_n517), .C1(new_n522), .C2(new_n521), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n605), .A2(G179), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT30), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n680), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT97), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT97), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n696), .B(new_n680), .C1(new_n687), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n579), .A2(new_n621), .A3(new_n658), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT31), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT98), .B1(new_n685), .B2(new_n686), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n687), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(KEYINPUT98), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n651), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n698), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT99), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT99), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n699), .A2(KEYINPUT31), .B1(new_n704), .B2(new_n651), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n709), .B(G330), .C1(new_n710), .C2(new_n698), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n678), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n676), .B1(new_n713), .B2(G1), .ZN(G364));
  INV_X1    g0514(.A(G13), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G45), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT101), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(KEYINPUT101), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n671), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n670), .A2(new_n325), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT102), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n724), .A2(G355), .B1(new_n515), .B2(new_n670), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n233), .A2(new_n485), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n670), .A2(new_n265), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(new_n485), .C2(new_n248), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n277), .B1(new_n212), .B2(G169), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT103), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT103), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n722), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n733), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n212), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n423), .A3(G200), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G107), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n212), .A2(new_n349), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n423), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G50), .A2(new_n749), .B1(new_n751), .B2(G68), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n746), .B(new_n752), .C1(new_n220), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n423), .A2(G200), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT104), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n212), .A2(new_n349), .A3(KEYINPUT104), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n201), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n740), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G159), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n265), .B1(new_n765), .B2(KEYINPUT32), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n755), .A2(new_n349), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G97), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT32), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n764), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n754), .A2(new_n760), .A3(new_n766), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n761), .B1(new_n757), .B2(new_n758), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT105), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT105), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G77), .ZN(new_n778));
  INV_X1    g0578(.A(new_n762), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n779), .A2(G329), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n265), .B(new_n780), .C1(G326), .C2(new_n749), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n753), .B(KEYINPUT107), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G303), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n745), .A2(G283), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n768), .A2(G294), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n781), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G311), .B2(new_n777), .ZN(new_n787));
  INV_X1    g0587(.A(new_n759), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n788), .A2(G322), .B1(new_n751), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT108), .Z(new_n791));
  AOI22_X1  g0591(.A1(new_n772), .A2(new_n778), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n736), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n738), .B1(new_n739), .B2(new_n792), .C1(new_n654), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n654), .A2(G330), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT100), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n655), .A2(new_n722), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G396));
  NOR2_X1   g0598(.A1(new_n733), .A2(new_n734), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n722), .B1(new_n799), .B2(new_n364), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G137), .A2(new_n749), .B1(new_n751), .B2(G150), .ZN(new_n801));
  INV_X1    g0601(.A(G143), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n759), .C1(new_n776), .C2(new_n763), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n782), .A2(G50), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n745), .A2(G68), .ZN(new_n806));
  INV_X1    g0606(.A(G132), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n265), .B1(new_n762), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G58), .B2(new_n768), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G283), .A2(new_n751), .B1(new_n749), .B2(G303), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n265), .B1(new_n779), .B2(G311), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n811), .A2(new_n769), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G294), .B2(new_n788), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n744), .A2(new_n220), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G107), .B2(new_n782), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(new_n515), .C2(new_n776), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n629), .A2(new_n440), .A3(new_n651), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n440), .A2(new_n651), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n451), .A2(new_n456), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n800), .B1(new_n739), .B2(new_n818), .C1(new_n822), .C2(new_n735), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n708), .A2(new_n711), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n677), .A2(new_n819), .A3(new_n821), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n822), .A2(new_n643), .A3(new_n658), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n722), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n824), .A2(new_n827), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(G384));
  OAI21_X1  g0631(.A(new_n467), .B1(new_n464), .B2(new_n468), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT35), .ZN(new_n833));
  OAI211_X1 g0633(.A(G116), .B(new_n231), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  NAND3_X1  g0636(.A1(new_n232), .A2(G77), .A3(new_n302), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n838), .A2(KEYINPUT109), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(KEYINPUT109), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n207), .A2(G68), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT110), .Z(new_n842));
  NOR3_X1   g0642(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n715), .A2(G1), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n380), .A2(new_n651), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n403), .A2(new_n406), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n845), .B1(new_n403), .B2(new_n406), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n822), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n705), .A2(new_n679), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n710), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT40), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n649), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n347), .A2(new_n348), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n336), .A2(new_n337), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n342), .A2(KEYINPUT17), .A3(new_n292), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n625), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n339), .B(new_n291), .C1(new_n340), .C2(new_n341), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n856), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n623), .A2(new_n863), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n868), .B2(KEYINPUT113), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT113), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n870), .B(new_n866), .C1(new_n856), .C2(new_n867), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n861), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n333), .A2(new_n316), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n263), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT112), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(KEYINPUT112), .A3(new_n263), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n855), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n362), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n352), .A3(new_n879), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n880), .A3(new_n336), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n865), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n874), .A2(new_n887), .ZN(new_n888));
  AOI221_X4 g0688(.A(new_n873), .B1(new_n865), .B2(new_n885), .C1(new_n362), .C2(new_n881), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n882), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n852), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(KEYINPUT114), .B(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n854), .A2(new_n888), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n851), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n458), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(G330), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n894), .B1(new_n458), .B2(new_n895), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n336), .B1(new_n342), .B2(new_n351), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n359), .A2(new_n360), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n855), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n870), .B1(new_n903), .B2(new_n866), .ZN(new_n904));
  OAI211_X1 g0704(.A(KEYINPUT113), .B(KEYINPUT37), .C1(new_n857), .C2(new_n901), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n865), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n906), .B2(new_n861), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n900), .B1(new_n907), .B2(new_n889), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n627), .A2(new_n380), .A3(new_n658), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n890), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n456), .A2(new_n651), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT111), .Z(new_n915));
  NAND2_X1  g0715(.A1(new_n826), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n847), .A2(new_n848), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n911), .A2(new_n887), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n625), .B2(new_n649), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n678), .A2(new_n458), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n636), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n899), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n211), .B2(new_n716), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n899), .A2(new_n926), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n836), .B1(new_n843), .B2(new_n844), .C1(new_n928), .C2(new_n929), .ZN(G367));
  NAND2_X1  g0730(.A1(new_n478), .A2(new_n651), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n502), .A2(new_n538), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n502), .B2(new_n658), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n667), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT44), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n667), .A2(new_n934), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n663), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n662), .A2(new_n664), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n666), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n655), .B(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n713), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT117), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n678), .A2(new_n712), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT117), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n713), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n671), .B(KEYINPUT41), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n720), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n666), .A2(new_n934), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n502), .B1(new_n932), .B2(new_n657), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n957), .A2(new_n958), .B1(new_n658), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n525), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n528), .A2(new_n658), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT115), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n639), .C2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n963), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n960), .A2(KEYINPUT116), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT116), .B1(new_n960), .B2(new_n968), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n966), .B(new_n967), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n969), .A2(new_n970), .B1(new_n960), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n940), .A2(new_n934), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n972), .B(new_n973), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n955), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n727), .A2(new_n241), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n737), .B1(new_n215), .B2(new_n435), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n745), .A2(G97), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n782), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n325), .B1(new_n762), .B2(new_n982), .C1(new_n750), .C2(new_n559), .ZN(new_n983));
  INV_X1    g0783(.A(new_n768), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(new_n446), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(G311), .C2(new_n749), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n753), .A2(new_n515), .ZN(new_n987));
  INV_X1    g0787(.A(G303), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n986), .B1(KEYINPUT46), .B2(new_n987), .C1(new_n988), .C2(new_n759), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n981), .B(new_n989), .C1(G283), .C2(new_n777), .ZN(new_n990));
  INV_X1    g0790(.A(G137), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n265), .B1(new_n762), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n984), .A2(new_n202), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n788), .C2(G150), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n748), .A2(new_n802), .B1(new_n753), .B2(new_n201), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G159), .B2(new_n751), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(new_n364), .C2(new_n744), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G50), .B2(new_n777), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n990), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT47), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n733), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(KEYINPUT47), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n721), .B1(new_n977), .B2(new_n978), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT118), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n966), .A2(new_n736), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n976), .A2(new_n1007), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n948), .A2(new_n950), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n671), .C1(new_n713), .C2(new_n945), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n720), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n793), .B1(new_n660), .B2(new_n661), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n777), .A2(G68), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n768), .A2(new_n434), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n265), .C1(new_n409), .C2(new_n762), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n753), .A2(new_n364), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n763), .B2(new_n748), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n788), .A2(G50), .B1(new_n251), .B2(new_n751), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1013), .A2(new_n979), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n265), .B1(new_n779), .B2(G326), .ZN(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n984), .A2(new_n1022), .B1(new_n559), .B2(new_n753), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G311), .A2(new_n751), .B1(new_n749), .B2(G322), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n982), .B2(new_n759), .C1(new_n776), .C2(new_n988), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1021), .B1(new_n515), .B2(new_n744), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n733), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n737), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n727), .B1(new_n238), .B2(new_n485), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n724), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n674), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n250), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT50), .B1(new_n250), .B2(G50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n674), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1037), .A2(new_n1041), .B1(new_n446), .B2(new_n670), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1033), .B(new_n721), .C1(new_n1034), .C2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1010), .B1(new_n1011), .B2(new_n944), .C1(new_n1012), .C2(new_n1043), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n951), .A2(new_n671), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n941), .B1(new_n950), .B2(new_n948), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n934), .A2(new_n736), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n737), .B1(new_n384), .B2(new_n215), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n727), .A2(new_n245), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n721), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n265), .B1(new_n762), .B2(new_n802), .C1(new_n202), .C2(new_n753), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n768), .A2(G77), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n207), .B2(new_n750), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n815), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n788), .A2(G159), .B1(G150), .B2(new_n749), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n776), .A2(new_n250), .B1(new_n1057), .B2(KEYINPUT51), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n788), .A2(G311), .B1(G317), .B2(new_n749), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT119), .B(KEYINPUT52), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n753), .A2(new_n1022), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n265), .B(new_n1064), .C1(G322), .C2(new_n779), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n751), .A2(G303), .B1(new_n768), .B2(G116), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n746), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n776), .A2(new_n559), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1059), .A2(new_n1060), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1052), .B1(new_n1069), .B2(new_n733), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n941), .A2(new_n720), .B1(new_n1049), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1047), .A2(new_n1048), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1048), .B1(new_n1047), .B2(new_n1071), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  NAND4_X1  g0876(.A1(new_n895), .A2(new_n918), .A3(G330), .A4(new_n822), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n910), .B1(new_n916), .B2(new_n918), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n908), .B2(new_n912), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n888), .A2(new_n1079), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1079), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT39), .B1(new_n874), .B2(new_n887), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n889), .A2(new_n890), .A3(new_n900), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n888), .A2(new_n1079), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n712), .A2(new_n822), .A3(new_n918), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n458), .A2(G330), .A3(new_n895), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n924), .A2(new_n636), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n918), .B1(new_n712), .B2(new_n822), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n916), .B1(new_n1093), .B2(new_n1078), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n895), .A2(G330), .A3(new_n822), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n919), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1088), .A2(new_n1096), .A3(new_n917), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1092), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1090), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1082), .A2(new_n1089), .A3(new_n1098), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n671), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n734), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n799), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n721), .B1(new_n1105), .B2(new_n251), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT121), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G107), .A2(new_n751), .B1(new_n749), .B2(G283), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n265), .B1(new_n779), .B2(G294), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1054), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n788), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n745), .A2(G68), .B1(new_n782), .B2(G87), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n384), .C2(new_n776), .ZN(new_n1113));
  INV_X1    g0913(.A(G125), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n265), .B1(new_n762), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G128), .B2(new_n749), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n763), .B2(new_n984), .C1(new_n744), .C2(new_n207), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n753), .A2(KEYINPUT53), .A3(new_n409), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT53), .B1(new_n753), .B2(new_n409), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n759), .B2(new_n807), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n776), .A2(new_n1122), .B1(new_n991), .B2(new_n750), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1124), .B2(KEYINPUT122), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT122), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1113), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1107), .B1(new_n1128), .B2(new_n733), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1103), .A2(new_n720), .B1(new_n1104), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1102), .A2(new_n1130), .ZN(G378));
  NAND2_X1  g0931(.A1(new_n415), .A2(new_n855), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n433), .B(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n894), .B2(G330), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n891), .A2(new_n893), .ZN(new_n1137));
  OAI211_X1 g0937(.A(KEYINPUT40), .B(new_n852), .C1(new_n907), .C2(new_n889), .ZN(new_n1138));
  AND4_X1   g0938(.A1(G330), .A2(new_n1137), .A3(new_n1138), .A4(new_n1135), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n923), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n913), .A2(new_n922), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1137), .A2(new_n1138), .A3(G330), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1135), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n894), .A2(G330), .A3(new_n1135), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1092), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1101), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n1149), .A3(KEYINPUT57), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n671), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT57), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n748), .A2(new_n1114), .B1(new_n753), .B2(new_n1122), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n984), .A2(new_n409), .B1(new_n807), .B2(new_n750), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G128), .C2(new_n788), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n991), .B2(new_n776), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT59), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1158), .A2(KEYINPUT123), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(KEYINPUT123), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n779), .C2(G124), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n744), .B2(new_n763), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n265), .A2(G41), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1164), .B1(new_n1022), .B2(new_n762), .C1(new_n984), .C2(new_n202), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1016), .B1(new_n384), .B2(new_n750), .C1(new_n515), .C2(new_n748), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(G107), .C2(new_n788), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n201), .B2(new_n744), .C1(new_n435), .C2(new_n776), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n733), .B1(new_n1163), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT124), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n722), .B1(new_n799), .B2(new_n207), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n1135), .C2(new_n735), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT125), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1147), .B2(new_n720), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1153), .A2(new_n1180), .ZN(G375));
  NAND3_X1  g0981(.A1(new_n1094), .A2(new_n1092), .A3(new_n1097), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1099), .A2(new_n954), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n919), .A2(new_n734), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n721), .B1(new_n1105), .B2(G68), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G116), .A2(new_n751), .B1(new_n749), .B2(G294), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n265), .B1(new_n779), .B2(G303), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1014), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G283), .B2(new_n788), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n745), .A2(G77), .B1(new_n782), .B2(G97), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n446), .C2(new_n776), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n776), .A2(new_n409), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n745), .A2(G58), .B1(new_n782), .B2(G159), .ZN(new_n1194));
  INV_X1    g0994(.A(G128), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n265), .B1(new_n762), .B2(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n807), .A2(new_n748), .B1(new_n750), .B2(new_n1122), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G50), .C2(new_n768), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1194), .B(new_n1198), .C1(new_n991), .C2(new_n759), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1192), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1186), .B1(new_n1200), .B2(new_n733), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1184), .A2(new_n720), .B1(new_n1185), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1183), .A2(new_n1202), .ZN(G381));
  OR2_X1    g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(G387), .A2(new_n1204), .A3(G384), .A4(G381), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1102), .A2(new_n1130), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1075), .A3(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(G375), .ZN(G407));
  NAND2_X1  g1008(.A1(new_n650), .A2(G213), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G407), .B(G213), .C1(G375), .C2(new_n1211), .ZN(G409));
  INV_X1    g1012(.A(new_n1074), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(G387), .A2(new_n1072), .A3(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(G393), .B(G396), .Z(new_n1215));
  OAI211_X1 g1015(.A(new_n976), .B(new_n1007), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1215), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT63), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G378), .B(new_n1180), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1147), .A2(new_n1149), .A3(new_n954), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1147), .A2(new_n720), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1178), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1206), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1209), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G384), .B(KEYINPUT126), .Z(new_n1228));
  INV_X1    g1028(.A(KEYINPUT60), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1184), .A2(new_n1229), .A3(new_n1148), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1230), .A2(G41), .A3(new_n670), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1182), .B1(new_n1098), .B2(new_n1229), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1228), .B1(new_n1233), .B2(new_n1202), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1202), .ZN(new_n1235));
  OR2_X1    g1035(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1235), .B(new_n1237), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1220), .B1(new_n1227), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1210), .A2(G2897), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(new_n1202), .A3(new_n1236), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1235), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1242), .C1(new_n1246), .C2(new_n1228), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1227), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1210), .B1(new_n1221), .B2(new_n1225), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1239), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1219), .A2(new_n1241), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1250), .A2(new_n1253), .A3(new_n1239), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1250), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1250), .B2(new_n1239), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1254), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1252), .B1(new_n1259), .B2(new_n1219), .ZN(G405));
  AOI21_X1  g1060(.A(G378), .B1(new_n1153), .B2(new_n1180), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1221), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1239), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1239), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1264), .A2(new_n1265), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1219), .A3(new_n1263), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(G402));
endmodule


