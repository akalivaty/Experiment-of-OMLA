//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(G1gat), .ZN(new_n205));
  AOI21_X1  g004(.A(G8gat), .B1(new_n205), .B2(KEYINPUT96), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n206), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G43gat), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n224));
  OAI21_X1  g023(.A(G36gat), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n215), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n213), .A2(G50gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n211), .A2(G43gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n230), .A2(new_n225), .A3(new_n215), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n218), .A2(new_n220), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT94), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT94), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n210), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n228), .A2(new_n229), .A3(new_n227), .ZN(new_n240));
  OR2_X1    g039(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n217), .B1(new_n241), .B2(new_n222), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(new_n242), .B2(new_n232), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT94), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT94), .B1(new_n218), .B2(new_n220), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n225), .A3(new_n215), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n248), .A2(KEYINPUT95), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT95), .B1(new_n248), .B2(new_n249), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n210), .B(new_n239), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT97), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n237), .B2(KEYINPUT17), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n248), .A2(KEYINPUT95), .A3(new_n249), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(KEYINPUT97), .A3(new_n210), .A4(new_n239), .ZN(new_n259));
  AOI211_X1 g058(.A(new_n203), .B(new_n238), .C1(new_n254), .C2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT99), .B1(new_n260), .B2(KEYINPUT18), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G141gat), .ZN(new_n262));
  INV_X1    g061(.A(G197gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT11), .B(G169gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n266), .B(KEYINPUT12), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n210), .B(new_n237), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n202), .B(KEYINPUT13), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n260), .B2(KEYINPUT18), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n259), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT18), .B(new_n202), .C1(new_n210), .C2(new_n237), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT98), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT98), .ZN(new_n276));
  AOI211_X1 g075(.A(new_n276), .B(new_n273), .C1(new_n254), .C2(new_n259), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n261), .B(new_n267), .C1(new_n271), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(KEYINPUT98), .A3(new_n274), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n238), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(new_n202), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT18), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n285), .A2(new_n286), .B1(new_n268), .B2(new_n269), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT99), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n285), .B2(new_n286), .ZN(new_n289));
  INV_X1    g088(.A(new_n267), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n283), .B(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n279), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  INV_X1    g094(.A(G211gat), .ZN(new_n296));
  INV_X1    g095(.A(G218gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(KEYINPUT22), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300));
  AND2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT76), .B(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT2), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(G148gat), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n314), .A3(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n307), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT2), .B1(new_n320), .B2(new_n311), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n324), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  XOR2_X1   g125(.A(G155gat), .B(G162gat), .Z(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n310), .B2(new_n315), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n322), .B1(new_n328), .B2(new_n307), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n294), .B(new_n304), .C1(new_n332), .C2(KEYINPUT29), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT77), .B1(new_n324), .B2(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n326), .A3(new_n330), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n299), .B(new_n300), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT72), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT86), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(G228gat), .A3(G233gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n303), .A2(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n324), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n333), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n336), .A2(new_n337), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT3), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(KEYINPUT85), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n329), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n345), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n344), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT87), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G22gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G78gat), .B(G106gat), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT84), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT31), .B(G50gat), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n357), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n366), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G15gat), .B(G43gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT69), .ZN(new_n375));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n375), .B(G134gat), .C1(new_n376), .C2(KEYINPUT1), .ZN(new_n377));
  INV_X1    g176(.A(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G113gat), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G120gat), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT1), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G134gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G127gat), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n377), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n374), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(G134gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n376), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n391));
  OAI21_X1  g190(.A(G127gat), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT70), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G169gat), .ZN(new_n396));
  INV_X1    g195(.A(G176gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n398), .A2(KEYINPUT26), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(KEYINPUT26), .ZN(new_n401));
  INV_X1    g200(.A(G183gat), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT68), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT27), .B(G183gat), .Z(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT65), .B(G190gat), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT28), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT65), .B(G190gat), .Z(new_n411));
  INV_X1    g210(.A(KEYINPUT28), .ZN(new_n412));
  OR3_X1    g211(.A1(new_n402), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT27), .B1(new_n402), .B2(KEYINPUT67), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n407), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n410), .A2(new_n415), .A3(new_n407), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n406), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT25), .ZN(new_n420));
  INV_X1    g219(.A(new_n399), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n398), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT64), .B(G176gat), .Z(new_n424));
  NOR2_X1   g223(.A1(new_n422), .A2(G169gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT24), .B1(new_n402), .B2(new_n403), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT24), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(G183gat), .A3(G190gat), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n428), .A2(new_n430), .B1(new_n402), .B2(new_n403), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n420), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n411), .A2(new_n402), .B1(new_n428), .B2(new_n430), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n420), .B1(new_n425), .B2(new_n397), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n423), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n430), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(G183gat), .B2(new_n409), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT66), .A3(new_n423), .A4(new_n435), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n395), .B1(new_n419), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n410), .A2(new_n415), .A3(new_n407), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n405), .B1(new_n443), .B2(new_n416), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n394), .A4(new_n388), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n373), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n448), .B1(new_n442), .B2(new_n446), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT71), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n456), .A3(KEYINPUT32), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n450), .B(KEYINPUT32), .C1(new_n451), .C2(new_n373), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n448), .A3(new_n446), .ZN(new_n461));
  XOR2_X1   g260(.A(new_n461), .B(KEYINPUT34), .Z(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n462), .A3(new_n459), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n370), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G8gat), .B(G36gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n444), .A2(new_n445), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n444), .A2(new_n445), .B1(new_n347), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n338), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n347), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n419), .B2(new_n441), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n444), .A2(new_n445), .A3(new_n472), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n303), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n471), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n475), .A2(new_n479), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(new_n470), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(KEYINPUT30), .B2(new_n480), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n329), .B1(new_n386), .B2(new_n387), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT81), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n388), .A2(new_n394), .A3(new_n329), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n495));
  OAI211_X1 g294(.A(new_n491), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n340), .A2(new_n392), .A3(new_n393), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n332), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n332), .B2(new_n497), .ZN(new_n503));
  INV_X1    g302(.A(new_n489), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n494), .A2(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n329), .A2(new_n386), .A3(new_n387), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n500), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT79), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n511), .B(new_n500), .C1(new_n504), .C2(new_n508), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(KEYINPUT5), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n502), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G1gat), .B(G29gat), .Z(new_n515));
  XNOR2_X1  g314(.A(G57gat), .B(G85gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AND4_X1   g319(.A1(KEYINPUT83), .A2(new_n514), .A3(KEYINPUT6), .A4(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n509), .B2(KEYINPUT79), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n512), .C1(new_n506), .C2(new_n503), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n519), .B1(new_n524), .B2(new_n502), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT83), .B1(new_n525), .B2(KEYINPUT6), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n519), .A3(new_n502), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT82), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(new_n530), .A3(new_n519), .A4(new_n502), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n525), .A2(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n488), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT35), .B1(new_n467), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n485), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT37), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n471), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT38), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n470), .B1(new_n485), .B2(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n303), .B1(new_n473), .B2(new_n474), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n477), .A2(new_n338), .A3(new_n478), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT37), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n542), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n480), .B(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n541), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n527), .A2(new_n552), .A3(new_n534), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n368), .A2(new_n369), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n499), .B1(new_n496), .B2(new_n498), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n504), .A2(new_n508), .A3(new_n500), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT39), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(KEYINPUT89), .A3(KEYINPUT39), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n519), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT40), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n514), .A2(new_n520), .ZN(new_n569));
  INV_X1    g368(.A(new_n567), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n562), .A2(new_n519), .A3(new_n570), .A4(new_n564), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n488), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n554), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n488), .ZN(new_n574));
  AOI211_X1 g373(.A(KEYINPUT6), .B(new_n525), .C1(new_n529), .C2(new_n531), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT6), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n525), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n574), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n464), .A2(KEYINPUT36), .A3(new_n465), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n458), .A2(new_n462), .A3(new_n459), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n462), .B1(new_n458), .B2(new_n459), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n581), .A2(new_n370), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n536), .B1(new_n573), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n584), .A2(new_n585), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(new_n369), .A3(new_n368), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT92), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n554), .B2(new_n591), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n293), .B1(new_n588), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(G57gat), .A2(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G57gat), .A2(G64gat), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G71gat), .B(G78gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT9), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(KEYINPUT100), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n602), .A3(new_n601), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n599), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G127gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n210), .B1(new_n613), .B2(new_n612), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n306), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n258), .A2(new_n239), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G99gat), .A2(G106gat), .ZN(new_n636));
  INV_X1    g435(.A(G85gat), .ZN(new_n637));
  INV_X1    g436(.A(G92gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(KEYINPUT8), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n640), .B(new_n641), .C1(new_n637), .C2(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(G85gat), .A3(G92gat), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(KEYINPUT101), .B2(KEYINPUT7), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n635), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n640), .A2(new_n641), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n649), .A2(G85gat), .A3(G92gat), .A4(new_n644), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n650), .A2(new_n634), .A3(new_n642), .A4(new_n639), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n633), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G190gat), .B(G218gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n654), .A2(new_n248), .B1(KEYINPUT41), .B2(new_n628), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n655), .B2(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n632), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n661), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n631), .A3(new_n659), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n627), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT106), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n612), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n652), .A2(new_n612), .A3(KEYINPUT104), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n608), .A2(new_n611), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(KEYINPUT105), .A3(new_n651), .A4(new_n648), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n652), .B2(new_n612), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n654), .A2(KEYINPUT10), .A3(new_n674), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n668), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n678), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n668), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G120gat), .B(G148gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT107), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n690), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n683), .A2(new_n685), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n666), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n597), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n527), .A2(new_n534), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g499(.A(KEYINPUT108), .B(KEYINPUT16), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G8gat), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n696), .A2(new_n488), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(G8gat), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n696), .B2(new_n488), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(KEYINPUT42), .B2(new_n703), .ZN(G1325gat));
  INV_X1    g506(.A(G15gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n696), .A2(new_n708), .A3(new_n591), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n586), .A2(new_n582), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n696), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(new_n708), .ZN(G1326gat));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n370), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n627), .ZN(new_n717));
  INV_X1    g516(.A(new_n694), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n665), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n597), .A2(new_n721), .ZN(new_n722));
  NOR4_X1   g521(.A1(new_n722), .A2(new_n697), .A3(new_n224), .A4(new_n223), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT45), .Z(new_n724));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  INV_X1    g524(.A(new_n665), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n589), .B1(new_n581), .B2(new_n592), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n553), .A2(new_n554), .A3(new_n572), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n710), .B1(new_n535), .B2(new_n554), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n467), .A2(new_n594), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n592), .A2(KEYINPUT92), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n725), .B(new_n726), .C1(new_n730), .C2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n587), .A2(new_n573), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n596), .A2(new_n738), .A3(new_n727), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n739), .A2(new_n725), .A3(KEYINPUT44), .A4(new_n726), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n719), .A2(new_n293), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n742), .A2(new_n697), .B1(new_n224), .B2(new_n223), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n724), .A2(new_n743), .ZN(G1328gat));
  NAND4_X1  g543(.A1(new_n597), .A2(new_n217), .A3(new_n488), .A4(new_n721), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT46), .Z(new_n746));
  OAI21_X1  g545(.A(G36gat), .B1(new_n742), .B2(new_n574), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1329gat));
  OAI21_X1  g551(.A(new_n213), .B1(new_n722), .B2(new_n466), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n711), .A2(G43gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n742), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g555(.A(new_n211), .B1(new_n722), .B2(new_n554), .ZN(new_n757));
  NAND2_X1  g556(.A1(KEYINPUT112), .A2(KEYINPUT48), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n370), .A2(G50gat), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(new_n758), .C1(new_n742), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT112), .A2(KEYINPUT48), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n760), .B(new_n761), .Z(G1331gat));
  NOR3_X1   g561(.A1(new_n666), .A2(new_n292), .A3(new_n718), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n739), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n698), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n488), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n764), .A2(new_n771), .A3(new_n591), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n764), .A2(new_n711), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n771), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n764), .A2(new_n370), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n292), .A2(new_n627), .A3(new_n718), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n737), .A2(new_n740), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780), .B2(new_n697), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n292), .A2(new_n627), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n726), .B(new_n782), .C1(new_n730), .C2(new_n734), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n739), .A2(KEYINPUT51), .A3(new_n726), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n698), .A2(new_n637), .A3(new_n694), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n781), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1336gat));
  OAI21_X1  g591(.A(G92gat), .B1(new_n780), .B2(new_n574), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n785), .A2(KEYINPUT115), .A3(new_n786), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n795), .A3(new_n784), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n488), .A2(new_n638), .A3(new_n694), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n793), .B(new_n801), .C1(new_n788), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n780), .B2(new_n710), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n466), .A2(G99gat), .A3(new_n718), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n788), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1338gat));
  NOR3_X1   g607(.A1(new_n554), .A2(G106gat), .A3(new_n718), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n796), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT117), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n812), .A3(new_n796), .A4(new_n809), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n737), .A2(new_n740), .A3(new_n370), .A4(new_n779), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT53), .B1(new_n787), .B2(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n815), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n815), .A3(KEYINPUT118), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n817), .A2(new_n823), .ZN(G1339gat));
  NAND2_X1  g623(.A1(new_n695), .A2(new_n293), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n283), .A2(new_n287), .A3(new_n290), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n202), .B1(new_n272), .B2(new_n284), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n268), .A2(new_n269), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n266), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT119), .B(new_n266), .C1(new_n828), .C2(new_n829), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n827), .A2(new_n832), .A3(new_n694), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n680), .A2(new_n668), .A3(new_n681), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n682), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n680), .A2(new_n681), .ZN(new_n840));
  INV_X1    g639(.A(new_n668), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n690), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n836), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n680), .A2(new_n668), .A3(new_n681), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n692), .B1(new_n682), .B2(new_n838), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(KEYINPUT55), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n693), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n279), .B2(new_n291), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT120), .B1(new_n835), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n849), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n292), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n834), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n855), .A3(new_n665), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n726), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n827), .A2(new_n832), .A3(new_n833), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n826), .B1(new_n861), .B2(new_n717), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n697), .A2(new_n488), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n467), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(G113gat), .A3(new_n292), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n862), .A2(new_n697), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n593), .A2(new_n595), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n488), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n380), .B1(new_n872), .B2(new_n293), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n868), .A2(new_n873), .ZN(G1340gat));
  NAND3_X1  g673(.A1(new_n867), .A2(G120gat), .A3(new_n694), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n378), .B1(new_n872), .B2(new_n718), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(G1341gat));
  XNOR2_X1  g676(.A(KEYINPUT69), .B(G127gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n717), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n869), .A2(new_n627), .A3(new_n871), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n867), .A2(new_n879), .B1(new_n880), .B2(new_n878), .ZN(G1342gat));
  NAND2_X1  g680(.A1(new_n867), .A2(new_n726), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G134gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n872), .A2(G134gat), .A3(new_n665), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n710), .A2(new_n370), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n488), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n293), .A2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n869), .A2(KEYINPUT123), .A3(new_n889), .A4(new_n891), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n308), .A2(new_n309), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n864), .A2(new_n710), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n627), .B1(new_n856), .B2(new_n860), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n370), .B1(new_n899), .B2(new_n826), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n726), .B1(new_n853), .B2(new_n834), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n717), .B1(new_n903), .B2(new_n859), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT122), .B(new_n717), .C1(new_n903), .C2(new_n859), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n825), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n554), .A2(new_n901), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n898), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n897), .B1(new_n911), .B2(new_n292), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT58), .B1(new_n895), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n911), .B2(new_n292), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n900), .A2(new_n901), .B1(new_n908), .B2(new_n909), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n916), .A2(KEYINPUT124), .A3(new_n293), .A4(new_n898), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n915), .A2(new_n917), .A3(new_n897), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n890), .B2(new_n892), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n913), .B1(new_n918), .B2(new_n920), .ZN(G1344gat));
  NAND2_X1  g720(.A1(new_n863), .A2(new_n909), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n904), .A2(new_n825), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n901), .B1(new_n923), .B2(new_n554), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n864), .A2(new_n710), .A3(new_n694), .ZN(new_n926));
  OAI211_X1 g725(.A(KEYINPUT59), .B(G148gat), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT59), .B1(new_n890), .B2(new_n718), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n312), .A3(new_n314), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n930), .A3(new_n694), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(G1345gat));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n717), .A3(new_n898), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n627), .A2(new_n306), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n933), .A2(new_n306), .B1(new_n890), .B2(new_n934), .ZN(G1346gat));
  NOR2_X1   g734(.A1(new_n665), .A2(new_n305), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n869), .A2(new_n726), .A3(new_n889), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n911), .A2(new_n936), .B1(new_n937), .B2(new_n305), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n698), .A2(new_n574), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n467), .B(new_n939), .C1(new_n899), .C2(new_n826), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n940), .A2(new_n396), .A3(new_n293), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n862), .A2(new_n698), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n870), .A2(new_n574), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n292), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n941), .B1(new_n946), .B2(new_n396), .ZN(G1348gat));
  OAI21_X1  g746(.A(new_n397), .B1(new_n944), .B2(new_n718), .ZN(new_n948));
  INV_X1    g747(.A(new_n940), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n424), .A3(new_n694), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(G1349gat));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n949), .A2(new_n957), .A3(new_n627), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT126), .B1(new_n940), .B2(new_n717), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(G183gat), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n717), .A2(new_n408), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n961), .ZN(new_n962));
  AOI211_X1 g761(.A(new_n955), .B(new_n956), .C1(new_n960), .C2(new_n962), .ZN(new_n963));
  AND4_X1   g762(.A1(new_n954), .A2(new_n960), .A3(new_n962), .A4(KEYINPUT60), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n411), .A3(new_n726), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n726), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(G190gat), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n967), .B2(G190gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(G1351gat));
  NOR2_X1   g771(.A1(new_n888), .A2(new_n574), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n942), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n292), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n939), .A2(new_n710), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n977), .B1(new_n922), .B2(new_n924), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n293), .A2(new_n263), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  INV_X1    g779(.A(G204gat), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n694), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(KEYINPUT62), .B1(new_n974), .B2(new_n982), .ZN(new_n983));
  OR3_X1    g782(.A1(new_n974), .A2(KEYINPUT62), .A3(new_n982), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n978), .A2(new_n694), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n981), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n975), .A2(new_n296), .A3(new_n627), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n978), .A2(new_n627), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n297), .A3(new_n726), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n978), .A2(new_n726), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(new_n993), .B2(new_n297), .ZN(G1355gat));
endmodule


