//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT28), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR3_X1    g008(.A1(new_n209), .A2(KEYINPUT65), .A3(KEYINPUT26), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT65), .B1(new_n209), .B2(KEYINPUT26), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n206), .A2(new_n207), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n203), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT24), .A3(new_n207), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n207), .A2(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT25), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n218), .B(KEYINPUT64), .Z(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  INV_X1    g026(.A(new_n224), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n217), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n215), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G226gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT73), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT70), .ZN(new_n236));
  NAND2_X1  g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT22), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G197gat), .A2(G204gat), .ZN(new_n240));
  AND2_X1   g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT71), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n236), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n231), .B(KEYINPUT72), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n234), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n247), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n246), .A2(new_n231), .B1(new_n230), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(new_n244), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  INV_X1    g052(.A(G64gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT30), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n259), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G141gat), .B(G148gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT2), .ZN(new_n265));
  XNOR2_X1  g064(.A(G155gat), .B(G162gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(KEYINPUT74), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT75), .B(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G155gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n264), .B1(new_n270), .B2(KEYINPUT2), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT76), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT76), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G120gat), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT66), .B(G120gat), .Z(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n276), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n276), .A2(G120gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT1), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n279), .A2(KEYINPUT67), .A3(new_n280), .A4(new_n281), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n284), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n267), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT76), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(new_n272), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n284), .A2(new_n287), .A3(new_n288), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT4), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n296), .A3(KEYINPUT81), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n289), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT4), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n304), .B(new_n292), .C1(new_n293), .C2(new_n272), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n305), .A3(new_n295), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n301), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n297), .A2(new_n300), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT82), .B1(new_n312), .B2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n295), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n298), .A2(KEYINPUT79), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n294), .A2(new_n317), .A3(new_n295), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n308), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n291), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n275), .A2(new_n289), .A3(KEYINPUT78), .A4(new_n290), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT77), .B(KEYINPUT4), .C1(new_n294), .C2(new_n295), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n306), .A2(new_n308), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n321), .A2(new_n330), .A3(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G1gat), .B(G29gat), .Z(new_n333));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n314), .A2(new_n331), .A3(new_n337), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n263), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n244), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n305), .B2(new_n245), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G228gat), .ZN(new_n348));
  INV_X1    g147(.A(G233gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n304), .B1(new_n244), .B2(KEYINPUT29), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n294), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n347), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n242), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n236), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n236), .B2(new_n354), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT3), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n275), .A2(new_n357), .ZN(new_n358));
  OAI22_X1  g157(.A1(new_n346), .A2(new_n358), .B1(new_n348), .B2(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT83), .B1(new_n360), .B2(G22gat), .ZN(new_n361));
  XOR2_X1   g160(.A(G78gat), .B(G106gat), .Z(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT31), .ZN(new_n363));
  INV_X1    g162(.A(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G22gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(new_n367), .A3(new_n359), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n360), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n370), .B(new_n367), .C1(KEYINPUT83), .C2(new_n365), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n360), .A2(G22gat), .A3(new_n365), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT84), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n369), .A2(new_n371), .A3(KEYINPUT84), .A4(new_n372), .ZN(new_n376));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n230), .A2(new_n295), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n230), .A2(new_n295), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n383), .B2(KEYINPUT33), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT32), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n386), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n380), .A3(new_n382), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n391));
  NOR2_X1   g190(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n381), .A2(new_n380), .A3(new_n382), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n385), .B(new_n383), .C1(KEYINPUT33), .C2(new_n379), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n387), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n400), .A3(KEYINPUT69), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT69), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n398), .C1(new_n399), .C2(new_n387), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n375), .A2(new_n376), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n344), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT86), .B1(new_n405), .B2(KEYINPUT35), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n343), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n342), .A2(new_n343), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n408), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT35), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n375), .A2(new_n376), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n400), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n263), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n405), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n407), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n342), .B2(new_n343), .ZN(new_n419));
  INV_X1    g218(.A(new_n409), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n261), .B1(new_n260), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT38), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n251), .A2(new_n244), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n234), .A2(new_n248), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT37), .B(new_n425), .C1(new_n426), .C2(new_n244), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n249), .A2(KEYINPUT37), .A3(new_n252), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n257), .B1(new_n249), .B2(new_n252), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n421), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n259), .B(new_n431), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n301), .A2(new_n306), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n320), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(KEYINPUT39), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n436), .B(KEYINPUT39), .C1(new_n320), .C2(new_n319), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(new_n337), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n439), .B2(KEYINPUT40), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n339), .C1(KEYINPUT40), .C2(new_n439), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n441), .A3(new_n413), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n414), .A2(KEYINPUT36), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n401), .A2(KEYINPUT36), .A3(new_n403), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n413), .B2(new_n344), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n418), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G22gat), .ZN(new_n451));
  INV_X1    g250(.A(G1gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT16), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n451), .A2(G1gat), .ZN(new_n455));
  OAI21_X1  g254(.A(G8gat), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n453), .ZN(new_n457));
  INV_X1    g256(.A(G8gat), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n457), .B(new_n458), .C1(G1gat), .C2(new_n451), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT9), .ZN(new_n461));
  INV_X1    g260(.A(G71gat), .ZN(new_n462));
  INV_X1    g261(.A(G78gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n254), .A2(G57gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n254), .A2(G57gat), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n464), .B(KEYINPUT93), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G78gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G57gat), .B(G64gat), .Z(new_n471));
  NAND4_X1  g270(.A1(new_n471), .A2(KEYINPUT93), .A3(new_n468), .A4(new_n464), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n460), .B1(KEYINPUT21), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G183gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(G231gat), .A2(G233gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G127gat), .B(G155gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(G211gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n478), .B(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n474), .A2(KEYINPUT21), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n482), .B(new_n483), .Z(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n481), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487));
  INV_X1    g286(.A(G29gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(G36gat), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G29gat), .B2(G36gat), .ZN(new_n493));
  INV_X1    g292(.A(G36gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n488), .A2(new_n494), .A3(KEYINPUT14), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT89), .B1(new_n500), .B2(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n497), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n502), .A2(new_n491), .A3(new_n493), .A4(new_n495), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n491), .A2(new_n495), .ZN(new_n505));
  INV_X1    g304(.A(new_n499), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n502), .A4(new_n493), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n256), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT8), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G99gat), .B(G106gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n513), .A2(new_n516), .A3(new_n520), .A4(new_n518), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n504), .A2(KEYINPUT17), .A3(new_n507), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(G99gat), .B2(G106gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(G85gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n256), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n520), .B1(new_n531), .B2(new_n513), .ZN(new_n532));
  INV_X1    g331(.A(new_n523), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n527), .B1(new_n508), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G190gat), .B(G218gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT95), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT96), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n536), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n539), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n536), .B2(new_n539), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n536), .A2(new_n539), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n524), .A2(new_n473), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n522), .A2(new_n523), .A3(new_n472), .A4(new_n470), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n556), .B2(new_n555), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n534), .A2(new_n474), .A3(KEYINPUT98), .A4(KEYINPUT10), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n554), .B2(new_n556), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT100), .B(G148gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(G120gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n564), .B1(new_n561), .B2(new_n562), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT101), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n574), .A2(new_n575), .A3(new_n571), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n574), .B2(new_n571), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n486), .A2(new_n553), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT102), .ZN(new_n581));
  INV_X1    g380(.A(new_n460), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n510), .A2(new_n525), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT90), .Z(new_n585));
  AOI21_X1  g384(.A(KEYINPUT91), .B1(new_n508), .B2(new_n460), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n508), .A2(KEYINPUT91), .A3(new_n460), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n583), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT92), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT18), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n587), .A2(new_n586), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n507), .A3(new_n504), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n585), .B(KEYINPUT13), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(KEYINPUT92), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n590), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n590), .A2(new_n596), .A3(new_n598), .A4(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n450), .A2(new_n581), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n410), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n263), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT16), .B(G8gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT103), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n615), .A2(KEYINPUT42), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(G8gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(KEYINPUT42), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(G1325gat));
  INV_X1    g418(.A(new_n414), .ZN(new_n620));
  AOI21_X1  g419(.A(G15gat), .B1(new_n610), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n445), .A2(G15gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT104), .Z(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n610), .B2(new_n623), .ZN(G1326gat));
  INV_X1    g423(.A(new_n413), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT43), .B(G22gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1327gat));
  AND2_X1   g427(.A1(new_n489), .A2(new_n490), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n412), .B(new_n415), .C1(new_n419), .C2(new_n420), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n625), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT86), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n633), .B(new_n412), .C1(new_n344), .C2(new_n404), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n632), .A2(new_n406), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n625), .B1(new_n421), .B2(new_n432), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n447), .B1(new_n636), .B2(new_n441), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n630), .B(new_n552), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n450), .A2(new_n630), .A3(KEYINPUT44), .A4(new_n552), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n609), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n486), .A2(new_n578), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n410), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n629), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n450), .A2(new_n552), .A3(new_n644), .ZN(new_n648));
  INV_X1    g447(.A(new_n629), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n410), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT45), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(G1328gat));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n494), .A3(new_n263), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT46), .Z(new_n654));
  OAI21_X1  g453(.A(G36gat), .B1(new_n645), .B2(new_n434), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(G1329gat));
  AND3_X1   g455(.A1(new_n648), .A2(new_n500), .A3(new_n620), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n445), .A3(new_n644), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n658), .B2(G43gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n660));
  OR2_X1    g459(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(G1330gat));
  NAND4_X1  g463(.A1(new_n640), .A2(new_n625), .A3(new_n641), .A4(new_n644), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n364), .B1(new_n665), .B2(KEYINPUT107), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(KEYINPUT107), .B2(new_n665), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n648), .A2(new_n364), .A3(new_n625), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT48), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(G50gat), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n670), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(KEYINPUT48), .B2(new_n671), .ZN(G1331gat));
  XNOR2_X1  g471(.A(new_n481), .B(new_n484), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n552), .ZN(new_n674));
  AND4_X1   g473(.A1(new_n674), .A2(new_n450), .A3(new_n578), .A4(new_n643), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n410), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT108), .B(G57gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1332gat));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n263), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT49), .B(G64gat), .Z(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(G1333gat));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n462), .A3(new_n620), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n675), .A2(new_n445), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n462), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g485(.A1(new_n675), .A2(new_n625), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n643), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT109), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n640), .A2(new_n578), .A3(new_n641), .A4(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n646), .A3(new_n530), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n553), .B(new_n690), .C1(new_n418), .C2(new_n449), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(KEYINPUT51), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(KEYINPUT51), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n579), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n410), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n693), .B1(new_n698), .B2(new_n530), .ZN(G1336gat));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n578), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n256), .B1(new_n701), .B2(new_n434), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n692), .A2(new_n256), .A3(new_n434), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(KEYINPUT52), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n706));
  AOI21_X1  g505(.A(G92gat), .B1(new_n697), .B2(new_n263), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n703), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1337gat));
  OAI21_X1  g508(.A(G99gat), .B1(new_n692), .B2(new_n446), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n701), .A2(G99gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n414), .ZN(G1338gat));
  OAI21_X1  g511(.A(G106gat), .B1(new_n692), .B2(new_n413), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT110), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n413), .A2(G106gat), .A3(new_n579), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT111), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n718), .B(G106gat), .C1(new_n692), .C2(new_n413), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT53), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n692), .A2(new_n722), .A3(new_n413), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n692), .B2(new_n413), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(G106gat), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n726), .A3(new_n717), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n727), .ZN(G1339gat));
  INV_X1    g527(.A(KEYINPUT118), .ZN(new_n729));
  INV_X1    g528(.A(new_n562), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n557), .A2(new_n560), .A3(new_n559), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n563), .A2(KEYINPUT54), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT54), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n561), .A2(new_n733), .A3(new_n562), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n734), .A2(KEYINPUT114), .A3(new_n572), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT114), .B1(new_n734), .B2(new_n572), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT55), .B(new_n732), .C1(new_n735), .C2(new_n736), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT101), .B1(new_n566), .B2(new_n572), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n574), .A2(new_n575), .A3(new_n571), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n740), .A2(new_n743), .A3(KEYINPUT115), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT115), .B1(new_n740), .B2(new_n743), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n609), .B(new_n739), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n585), .B1(new_n591), .B2(new_n583), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n592), .B(new_n594), .C1(new_n587), .C2(new_n586), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n604), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n608), .A2(new_n578), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT116), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n608), .A2(new_n578), .A3(new_n753), .A4(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n746), .A2(new_n755), .A3(KEYINPUT117), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n553), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n608), .A2(new_n750), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n761), .B(new_n739), .C1(new_n744), .C2(new_n745), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n553), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n486), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n580), .B2(new_n609), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n674), .A2(KEYINPUT113), .A3(new_n643), .A4(new_n579), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n729), .B1(new_n770), .B2(new_n625), .ZN(new_n771));
  OAI211_X1 g570(.A(KEYINPUT118), .B(new_n413), .C1(new_n765), .C2(new_n769), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n646), .A2(new_n263), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(new_n620), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G113gat), .B1(new_n775), .B2(new_n643), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n746), .A2(KEYINPUT117), .A3(new_n755), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT117), .B1(new_n746), .B2(new_n755), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(new_n552), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n673), .B1(new_n779), .B2(new_n763), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n767), .A2(new_n768), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n401), .A2(new_n403), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n413), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n774), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n276), .A3(new_n609), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n776), .A2(new_n788), .ZN(G1340gat));
  OAI21_X1  g588(.A(G120gat), .B1(new_n775), .B2(new_n579), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n579), .A2(new_n278), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n786), .B2(new_n791), .ZN(G1341gat));
  INV_X1    g591(.A(G127gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n775), .A2(new_n793), .A3(new_n673), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n786), .A2(new_n673), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT119), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n793), .ZN(G1342gat));
  NOR3_X1   g596(.A1(new_n786), .A2(G134gat), .A3(new_n553), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT120), .Z(new_n801));
  OAI21_X1  g600(.A(G134gat), .B1(new_n775), .B2(new_n553), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n801), .B(new_n802), .C1(new_n799), .C2(new_n798), .ZN(G1343gat));
  NOR2_X1   g602(.A1(new_n770), .A2(new_n413), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n785), .A2(new_n445), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(G141gat), .A3(new_n643), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n804), .B2(KEYINPUT57), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810));
  OAI211_X1 g609(.A(KEYINPUT121), .B(new_n810), .C1(new_n770), .C2(new_n413), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n609), .A2(new_n743), .A3(new_n739), .A4(new_n740), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n751), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n553), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n486), .B1(new_n764), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n625), .C1(new_n769), .C2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n809), .A2(new_n811), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n609), .A3(new_n805), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n807), .B1(new_n818), .B2(G141gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1344gat));
  NOR3_X1   g622(.A1(new_n806), .A2(G148gat), .A3(new_n579), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT123), .ZN(new_n825));
  INV_X1    g624(.A(G148gat), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n817), .A2(new_n805), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT59), .B(new_n826), .C1(new_n827), .C2(new_n578), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n581), .A2(new_n643), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n810), .B(new_n625), .C1(new_n830), .C2(new_n815), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT57), .B1(new_n770), .B2(new_n413), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n578), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n805), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(G148gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n825), .B1(new_n828), .B2(new_n836), .ZN(G1345gat));
  NAND3_X1  g636(.A1(new_n827), .A2(G155gat), .A3(new_n486), .ZN(new_n838));
  INV_X1    g637(.A(G155gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n806), .B2(new_n673), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(G1346gat));
  NAND3_X1  g640(.A1(new_n827), .A2(new_n269), .A3(new_n552), .ZN(new_n842));
  INV_X1    g641(.A(new_n269), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n806), .B2(new_n553), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(G1347gat));
  NOR2_X1   g644(.A1(new_n410), .A2(new_n434), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n784), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(G169gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n609), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n414), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n773), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n773), .B2(new_n852), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(new_n643), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n850), .B1(new_n856), .B2(new_n849), .ZN(G1348gat));
  AOI21_X1  g656(.A(G176gat), .B1(new_n848), .B2(new_n578), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n854), .A2(new_n855), .A3(new_n579), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(G176gat), .ZN(G1349gat));
  AND2_X1   g659(.A1(new_n486), .A2(new_n202), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT125), .B1(new_n848), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n854), .A2(new_n855), .A3(new_n673), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n220), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n203), .A3(new_n552), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n782), .B2(new_n413), .ZN(new_n867));
  INV_X1    g666(.A(new_n772), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n852), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT124), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n552), .A3(new_n853), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n871), .A2(new_n872), .A3(G190gat), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n871), .B2(G190gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n866), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT126), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n866), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1351gat));
  NOR2_X1   g678(.A1(new_n847), .A2(new_n445), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n833), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G197gat), .B1(new_n882), .B2(new_n643), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n804), .A2(new_n880), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(G197gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n643), .B2(new_n885), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n834), .A2(new_n880), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G204gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n884), .A2(G204gat), .A3(new_n579), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1353gat));
  OR3_X1    g691(.A1(new_n884), .A2(G211gat), .A3(new_n673), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n881), .A2(new_n486), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT63), .B1(new_n894), .B2(G211gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1354gat));
  OAI21_X1  g696(.A(G218gat), .B1(new_n882), .B2(new_n553), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n884), .A2(G218gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n553), .B2(new_n899), .ZN(G1355gat));
endmodule


