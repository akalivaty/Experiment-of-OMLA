

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745;

  NAND2_X4 U368 ( .A1(n369), .A2(n366), .ZN(n508) );
  AND2_X2 U369 ( .A1(n577), .A2(n576), .ZN(n390) );
  AND2_X2 U370 ( .A1(n552), .A2(n568), .ZN(n567) );
  AND2_X2 U371 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X2 U372 ( .A(n388), .B(KEYINPUT45), .ZN(n365) );
  INV_X4 U373 ( .A(G128), .ZN(n414) );
  NAND2_X1 U374 ( .A1(n409), .A2(n406), .ZN(n626) );
  AND2_X1 U375 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U376 ( .A(n392), .B(n391), .ZN(n744) );
  OR2_X1 U377 ( .A1(n672), .A2(n522), .ZN(n392) );
  XNOR2_X1 U378 ( .A(n396), .B(n395), .ZN(n660) );
  NOR2_X1 U379 ( .A1(n600), .A2(G902), .ZN(n467) );
  INV_X1 U380 ( .A(n379), .ZN(n345) );
  XNOR2_X1 U381 ( .A(n372), .B(n355), .ZN(n400) );
  BUF_X1 U382 ( .A(n360), .Z(n346) );
  NAND2_X1 U383 ( .A1(n365), .A2(n387), .ZN(n677) );
  XNOR2_X2 U384 ( .A(n467), .B(n374), .ZN(n581) );
  XNOR2_X2 U385 ( .A(n500), .B(n499), .ZN(n691) );
  NAND2_X1 U386 ( .A1(n527), .A2(n382), .ZN(n381) );
  NOR2_X1 U387 ( .A1(G953), .A2(G237), .ZN(n461) );
  XNOR2_X1 U388 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n417) );
  XNOR2_X1 U389 ( .A(n440), .B(n348), .ZN(n731) );
  OR2_X1 U390 ( .A1(n659), .A2(n553), .ZN(n554) );
  NOR2_X1 U391 ( .A1(n661), .A2(n354), .ZN(n405) );
  AND2_X1 U392 ( .A1(n526), .A2(n624), .ZN(n382) );
  INV_X1 U393 ( .A(G469), .ZN(n368) );
  NAND2_X1 U394 ( .A1(G902), .A2(G469), .ZN(n370) );
  XNOR2_X1 U395 ( .A(n465), .B(n463), .ZN(n378) );
  XOR2_X1 U396 ( .A(KEYINPUT79), .B(KEYINPUT93), .Z(n463) );
  XNOR2_X1 U397 ( .A(n462), .B(n464), .ZN(n377) );
  XNOR2_X1 U398 ( .A(G113), .B(G116), .ZN(n464) );
  NAND2_X1 U399 ( .A1(n519), .A2(n347), .ZN(n394) );
  NOR2_X1 U400 ( .A1(n744), .A2(n745), .ZN(n518) );
  XNOR2_X1 U401 ( .A(G140), .B(KEYINPUT11), .ZN(n418) );
  XOR2_X1 U402 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n419) );
  XNOR2_X1 U403 ( .A(n421), .B(n364), .ZN(n363) );
  INV_X1 U404 ( .A(KEYINPUT98), .ZN(n364) );
  XNOR2_X1 U405 ( .A(G131), .B(G143), .ZN(n421) );
  INV_X1 U406 ( .A(G137), .ZN(n398) );
  XNOR2_X1 U407 ( .A(n460), .B(G101), .ZN(n481) );
  XNOR2_X1 U408 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n460) );
  XNOR2_X1 U409 ( .A(G119), .B(KEYINPUT3), .ZN(n459) );
  XOR2_X1 U410 ( .A(G116), .B(G107), .Z(n486) );
  INV_X1 U411 ( .A(G472), .ZN(n374) );
  XNOR2_X1 U412 ( .A(n384), .B(n383), .ZN(n439) );
  INV_X1 U413 ( .A(KEYINPUT8), .ZN(n383) );
  XNOR2_X1 U414 ( .A(n506), .B(KEYINPUT41), .ZN(n672) );
  NOR2_X1 U415 ( .A1(n660), .A2(n659), .ZN(n506) );
  NAND2_X1 U416 ( .A1(n379), .A2(n412), .ZN(n410) );
  NOR2_X1 U417 ( .A1(n713), .A2(G902), .ZN(n445) );
  OR2_X1 U418 ( .A1(n708), .A2(G902), .ZN(n434) );
  XNOR2_X1 U419 ( .A(n427), .B(n362), .ZN(n528) );
  XNOR2_X1 U420 ( .A(n426), .B(G475), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n543), .B(KEYINPUT0), .ZN(n544) );
  BUF_X1 U422 ( .A(n581), .Z(n358) );
  XNOR2_X1 U423 ( .A(n581), .B(n373), .ZN(n588) );
  INV_X1 U424 ( .A(KEYINPUT6), .ZN(n373) );
  INV_X1 U425 ( .A(KEYINPUT77), .ZN(n413) );
  INV_X1 U426 ( .A(n661), .ZN(n524) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n448) );
  INV_X1 U428 ( .A(n581), .ZN(n646) );
  INV_X1 U429 ( .A(KEYINPUT105), .ZN(n395) );
  NAND2_X1 U430 ( .A1(n657), .A2(n656), .ZN(n396) );
  INV_X1 U431 ( .A(G237), .ZN(n469) );
  NAND2_X1 U432 ( .A1(n368), .A2(n470), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n466), .B(n376), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n394), .B(n393), .ZN(n386) );
  XNOR2_X1 U436 ( .A(n594), .B(n593), .ZN(n389) );
  XNOR2_X1 U437 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U438 ( .A(n420), .B(n363), .ZN(n424) );
  XNOR2_X1 U439 ( .A(n484), .B(n415), .ZN(n423) );
  XNOR2_X1 U440 ( .A(n497), .B(n397), .ZN(n499) );
  XNOR2_X1 U441 ( .A(n399), .B(n348), .ZN(n397) );
  XNOR2_X1 U442 ( .A(n498), .B(n496), .ZN(n399) );
  XNOR2_X1 U443 ( .A(n481), .B(n480), .ZN(n497) );
  XNOR2_X1 U444 ( .A(KEYINPUT73), .B(G110), .ZN(n480) );
  INV_X1 U445 ( .A(KEYINPUT80), .ZN(n510) );
  XNOR2_X1 U446 ( .A(n600), .B(KEYINPUT62), .ZN(n601) );
  XNOR2_X1 U447 ( .A(n731), .B(n401), .ZN(n713) );
  XNOR2_X1 U448 ( .A(n403), .B(n402), .ZN(n401) );
  NAND2_X1 U449 ( .A1(n439), .A2(G221), .ZN(n402) );
  XNOR2_X1 U450 ( .A(n432), .B(n385), .ZN(n708) );
  XNOR2_X1 U451 ( .A(n431), .B(n433), .ZN(n385) );
  NOR2_X1 U452 ( .A1(n733), .A2(G952), .ZN(n717) );
  BUF_X1 U453 ( .A(G953), .Z(n359) );
  INV_X1 U454 ( .A(KEYINPUT42), .ZN(n391) );
  INV_X1 U455 ( .A(KEYINPUT40), .ZN(n516) );
  XNOR2_X1 U456 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n579) );
  NAND2_X1 U457 ( .A1(n408), .A2(n407), .ZN(n406) );
  AND2_X1 U458 ( .A1(n590), .A2(n589), .ZN(n614) );
  AND2_X1 U459 ( .A1(n380), .A2(n636), .ZN(n347) );
  XOR2_X1 U460 ( .A(n398), .B(G140), .Z(n348) );
  XOR2_X1 U461 ( .A(G131), .B(G134), .Z(n349) );
  XOR2_X1 U462 ( .A(n437), .B(KEYINPUT92), .Z(n350) );
  INV_X1 U463 ( .A(G146), .ZN(n458) );
  OR2_X1 U464 ( .A1(n542), .A2(n541), .ZN(n351) );
  XOR2_X1 U465 ( .A(n536), .B(KEYINPUT43), .Z(n352) );
  XOR2_X1 U466 ( .A(n586), .B(KEYINPUT96), .Z(n353) );
  XOR2_X1 U467 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n354) );
  XNOR2_X1 U468 ( .A(n521), .B(KEYINPUT19), .ZN(n355) );
  INV_X1 U469 ( .A(KEYINPUT84), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n500), .B(n375), .ZN(n600) );
  INV_X1 U471 ( .A(n493), .ZN(n356) );
  OR2_X1 U472 ( .A1(n537), .A2(n531), .ZN(n624) );
  BUF_X1 U473 ( .A(n697), .Z(n711) );
  XNOR2_X1 U474 ( .A(n346), .B(n539), .ZN(n357) );
  XNOR2_X1 U475 ( .A(n360), .B(n539), .ZN(n673) );
  NAND2_X1 U476 ( .A1(n578), .A2(n588), .ZN(n360) );
  XNOR2_X1 U477 ( .A(n537), .B(KEYINPUT38), .ZN(n657) );
  OR2_X1 U478 ( .A1(n584), .A2(n554), .ZN(n556) );
  AND2_X2 U479 ( .A1(n557), .A2(n639), .ZN(n578) );
  XNOR2_X1 U480 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U481 ( .A(n478), .B(n479), .ZN(n482) );
  NAND2_X1 U482 ( .A1(n573), .A2(n361), .ZN(n577) );
  NAND2_X1 U483 ( .A1(n571), .A2(n572), .ZN(n361) );
  XNOR2_X2 U484 ( .A(n556), .B(n555), .ZN(n563) );
  AND2_X1 U485 ( .A1(n365), .A2(n733), .ZN(n722) );
  OR2_X1 U486 ( .A1(n691), .A2(n367), .ZN(n366) );
  NAND2_X1 U487 ( .A1(n691), .A2(G469), .ZN(n371) );
  XNOR2_X2 U488 ( .A(n508), .B(KEYINPUT1), .ZN(n557) );
  NAND2_X1 U489 ( .A1(n400), .A2(n351), .ZN(n545) );
  NOR2_X2 U490 ( .A1(n537), .A2(n520), .ZN(n372) );
  XNOR2_X2 U491 ( .A(n492), .B(n491), .ZN(n537) );
  XNOR2_X2 U492 ( .A(n730), .B(G146), .ZN(n500) );
  XNOR2_X2 U493 ( .A(n478), .B(n349), .ZN(n730) );
  XNOR2_X2 U494 ( .A(n457), .B(n456), .ZN(n478) );
  AND2_X1 U495 ( .A1(n345), .A2(KEYINPUT84), .ZN(n407) );
  INV_X1 U496 ( .A(n400), .ZN(n379) );
  XNOR2_X1 U497 ( .A(n381), .B(n532), .ZN(n380) );
  NAND2_X1 U498 ( .A1(n733), .A2(G234), .ZN(n384) );
  INV_X4 U499 ( .A(G953), .ZN(n733) );
  INV_X1 U500 ( .A(n732), .ZN(n387) );
  NAND2_X1 U501 ( .A1(n386), .A2(n538), .ZN(n732) );
  NAND2_X1 U502 ( .A1(n390), .A2(n389), .ZN(n388) );
  NOR2_X2 U503 ( .A1(n673), .A2(n584), .ZN(n546) );
  INV_X1 U504 ( .A(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U505 ( .A(n438), .B(n350), .ZN(n403) );
  XNOR2_X1 U506 ( .A(n404), .B(n413), .ZN(n527) );
  NAND2_X1 U507 ( .A1(n626), .A2(n405), .ZN(n404) );
  INV_X1 U508 ( .A(n522), .ZN(n408) );
  NAND2_X1 U509 ( .A1(n522), .A2(n412), .ZN(n411) );
  XNOR2_X2 U510 ( .A(n414), .B(G143), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n704), .B(n703), .ZN(n706) );
  AND2_X2 U512 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X2 U513 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n474) );
  AND2_X1 U514 ( .A1(G214), .A2(n461), .ZN(n415) );
  AND2_X1 U515 ( .A1(n644), .A2(n454), .ZN(n416) );
  INV_X1 U516 ( .A(KEYINPUT76), .ZN(n532) );
  NOR2_X1 U517 ( .A1(n632), .A2(n617), .ZN(n586) );
  INV_X1 U518 ( .A(n614), .ZN(n591) );
  INV_X1 U519 ( .A(KEYINPUT24), .ZN(n437) );
  AND2_X1 U520 ( .A1(n564), .A2(n416), .ZN(n455) );
  NOR2_X1 U521 ( .A1(n582), .A2(n509), .ZN(n511) );
  XNOR2_X1 U522 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U523 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U524 ( .A(n517), .B(n516), .ZN(n745) );
  XNOR2_X1 U525 ( .A(n458), .B(G125), .ZN(n476) );
  XNOR2_X1 U526 ( .A(n476), .B(n417), .ZN(n440) );
  XNOR2_X1 U527 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U528 ( .A(G113), .B(G104), .ZN(n422) );
  XNOR2_X1 U529 ( .A(n422), .B(G122), .ZN(n484) );
  XNOR2_X1 U530 ( .A(n440), .B(n425), .ZN(n700) );
  NOR2_X1 U531 ( .A1(G902), .A2(n700), .ZN(n427) );
  XNOR2_X1 U532 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n426) );
  XNOR2_X1 U533 ( .A(n486), .B(KEYINPUT7), .ZN(n433) );
  XOR2_X1 U534 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n429) );
  NAND2_X1 U535 ( .A1(G217), .A2(n439), .ZN(n428) );
  XNOR2_X1 U536 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U537 ( .A(n430), .B(G122), .Z(n432) );
  XNOR2_X1 U538 ( .A(n457), .B(G134), .ZN(n431) );
  XNOR2_X1 U539 ( .A(G478), .B(n434), .ZN(n523) );
  NOR2_X1 U540 ( .A1(n528), .A2(n523), .ZN(n628) );
  INV_X1 U541 ( .A(n628), .ZN(n473) );
  XOR2_X1 U542 ( .A(KEYINPUT23), .B(G110), .Z(n436) );
  XNOR2_X1 U543 ( .A(G128), .B(G119), .ZN(n435) );
  XNOR2_X1 U544 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U545 ( .A(KEYINPUT25), .B(KEYINPUT81), .Z(n443) );
  XNOR2_X1 U546 ( .A(KEYINPUT15), .B(G902), .ZN(n595) );
  NAND2_X1 U547 ( .A1(G234), .A2(n595), .ZN(n441) );
  XNOR2_X1 U548 ( .A(KEYINPUT20), .B(n441), .ZN(n446) );
  NAND2_X1 U549 ( .A1(n446), .A2(G217), .ZN(n442) );
  XOR2_X1 U550 ( .A(n443), .B(n442), .Z(n444) );
  XNOR2_X2 U551 ( .A(n445), .B(n444), .ZN(n564) );
  AND2_X1 U552 ( .A1(n446), .A2(G221), .ZN(n447) );
  XNOR2_X1 U553 ( .A(n447), .B(KEYINPUT21), .ZN(n644) );
  XNOR2_X1 U554 ( .A(n448), .B(KEYINPUT14), .ZN(n449) );
  XNOR2_X1 U555 ( .A(KEYINPUT78), .B(n449), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n451), .A2(G952), .ZN(n450) );
  XOR2_X1 U557 ( .A(KEYINPUT91), .B(n450), .Z(n670) );
  NOR2_X1 U558 ( .A1(n670), .A2(n359), .ZN(n542) );
  AND2_X1 U559 ( .A1(n451), .A2(n359), .ZN(n452) );
  NAND2_X1 U560 ( .A1(G902), .A2(n452), .ZN(n540) );
  NOR2_X1 U561 ( .A1(G900), .A2(n540), .ZN(n453) );
  NOR2_X1 U562 ( .A1(n542), .A2(n453), .ZN(n509) );
  INV_X1 U563 ( .A(n509), .ZN(n454) );
  XNOR2_X1 U564 ( .A(n455), .B(KEYINPUT71), .ZN(n502) );
  INV_X1 U565 ( .A(KEYINPUT4), .ZN(n456) );
  XNOR2_X1 U566 ( .A(n459), .B(KEYINPUT72), .ZN(n483) );
  XNOR2_X1 U567 ( .A(n483), .B(n481), .ZN(n466) );
  NAND2_X1 U568 ( .A1(n461), .A2(G210), .ZN(n462) );
  XOR2_X1 U569 ( .A(G137), .B(KEYINPUT5), .Z(n465) );
  INV_X1 U570 ( .A(n588), .ZN(n468) );
  NOR2_X1 U571 ( .A1(n502), .A2(n468), .ZN(n471) );
  INV_X1 U572 ( .A(G902), .ZN(n470) );
  NAND2_X1 U573 ( .A1(n470), .A2(n469), .ZN(n490) );
  NAND2_X1 U574 ( .A1(n490), .A2(G214), .ZN(n656) );
  NAND2_X1 U575 ( .A1(n471), .A2(n656), .ZN(n472) );
  NOR2_X1 U576 ( .A1(n473), .A2(n472), .ZN(n534) );
  NAND2_X1 U577 ( .A1(n733), .A2(G224), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n482), .B(n497), .ZN(n489) );
  XNOR2_X1 U580 ( .A(n484), .B(n483), .ZN(n488) );
  INV_X1 U581 ( .A(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U582 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U583 ( .A(n488), .B(n487), .ZN(n723) );
  XNOR2_X1 U584 ( .A(n489), .B(n723), .ZN(n609) );
  NAND2_X1 U585 ( .A1(n609), .A2(n595), .ZN(n492) );
  NAND2_X1 U586 ( .A1(n490), .A2(G210), .ZN(n491) );
  INV_X1 U587 ( .A(n537), .ZN(n493) );
  NAND2_X1 U588 ( .A1(n534), .A2(n493), .ZN(n495) );
  XOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT36), .Z(n494) );
  XNOR2_X1 U590 ( .A(n495), .B(n494), .ZN(n501) );
  XNOR2_X1 U591 ( .A(G104), .B(G107), .ZN(n498) );
  NAND2_X1 U592 ( .A1(G227), .A2(n733), .ZN(n496) );
  NAND2_X1 U593 ( .A1(n501), .A2(n557), .ZN(n636) );
  NOR2_X1 U594 ( .A1(n502), .A2(n646), .ZN(n503) );
  XNOR2_X1 U595 ( .A(n503), .B(KEYINPUT28), .ZN(n505) );
  XNOR2_X1 U596 ( .A(n508), .B(KEYINPUT104), .ZN(n504) );
  NAND2_X1 U597 ( .A1(n505), .A2(n504), .ZN(n522) );
  INV_X1 U598 ( .A(n523), .ZN(n529) );
  NAND2_X1 U599 ( .A1(n528), .A2(n529), .ZN(n659) );
  NAND2_X1 U600 ( .A1(n581), .A2(n656), .ZN(n507) );
  XNOR2_X1 U601 ( .A(KEYINPUT30), .B(n507), .ZN(n513) );
  INV_X1 U602 ( .A(n644), .ZN(n553) );
  NOR2_X2 U603 ( .A1(n553), .A2(n564), .ZN(n639) );
  NAND2_X1 U604 ( .A1(n639), .A2(n508), .ZN(n582) );
  XNOR2_X1 U605 ( .A(n511), .B(n510), .ZN(n512) );
  NOR2_X1 U606 ( .A1(n513), .A2(n512), .ZN(n530) );
  AND2_X1 U607 ( .A1(n530), .A2(n657), .ZN(n515) );
  XNOR2_X1 U608 ( .A(KEYINPUT39), .B(KEYINPUT75), .ZN(n514) );
  XNOR2_X1 U609 ( .A(n515), .B(n514), .ZN(n533) );
  NAND2_X1 U610 ( .A1(n533), .A2(n628), .ZN(n517) );
  XNOR2_X1 U611 ( .A(n518), .B(KEYINPUT46), .ZN(n519) );
  INV_X1 U612 ( .A(n656), .ZN(n520) );
  INV_X1 U613 ( .A(KEYINPUT66), .ZN(n521) );
  AND2_X1 U614 ( .A1(n528), .A2(n523), .ZN(n631) );
  NOR2_X1 U615 ( .A1(n628), .A2(n631), .ZN(n661) );
  NAND2_X1 U616 ( .A1(n626), .A2(n524), .ZN(n525) );
  NAND2_X1 U617 ( .A1(n525), .A2(KEYINPUT47), .ZN(n526) );
  NOR2_X1 U618 ( .A1(n529), .A2(n528), .ZN(n547) );
  NAND2_X1 U619 ( .A1(n530), .A2(n547), .ZN(n531) );
  NAND2_X1 U620 ( .A1(n533), .A2(n631), .ZN(n637) );
  XNOR2_X1 U621 ( .A(KEYINPUT103), .B(n534), .ZN(n535) );
  NOR2_X1 U622 ( .A1(n557), .A2(n535), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n352), .A2(n356), .ZN(n607) );
  AND2_X1 U624 ( .A1(n637), .A2(n607), .ZN(n538) );
  XOR2_X1 U625 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n539) );
  NOR2_X1 U626 ( .A1(n540), .A2(G898), .ZN(n541) );
  INV_X1 U627 ( .A(KEYINPUT89), .ZN(n543) );
  XNOR2_X2 U628 ( .A(n545), .B(n544), .ZN(n584) );
  XNOR2_X1 U629 ( .A(n546), .B(KEYINPUT34), .ZN(n548) );
  NAND2_X1 U630 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X2 U631 ( .A(n549), .B(KEYINPUT35), .ZN(n743) );
  INV_X1 U632 ( .A(n743), .ZN(n551) );
  INV_X1 U633 ( .A(KEYINPUT88), .ZN(n550) );
  NAND2_X1 U634 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U635 ( .A(KEYINPUT44), .ZN(n568) );
  INV_X1 U636 ( .A(KEYINPUT22), .ZN(n555) );
  XNOR2_X1 U637 ( .A(n588), .B(KEYINPUT83), .ZN(n559) );
  XNOR2_X1 U638 ( .A(n564), .B(KEYINPUT101), .ZN(n643) );
  INV_X1 U639 ( .A(n557), .ZN(n641) );
  NOR2_X1 U640 ( .A1(n643), .A2(n641), .ZN(n558) );
  AND2_X1 U641 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U642 ( .A1(n563), .A2(n560), .ZN(n562) );
  XNOR2_X1 U643 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n561) );
  XNOR2_X1 U644 ( .A(n562), .B(n561), .ZN(n606) );
  AND2_X1 U645 ( .A1(n563), .A2(n641), .ZN(n590) );
  INV_X1 U646 ( .A(n564), .ZN(n565) );
  NOR2_X1 U647 ( .A1(n565), .A2(n358), .ZN(n566) );
  NAND2_X1 U648 ( .A1(n590), .A2(n566), .ZN(n621) );
  NAND2_X1 U649 ( .A1(n606), .A2(n621), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n567), .A2(n570), .ZN(n573) );
  NAND2_X1 U651 ( .A1(n568), .A2(KEYINPUT88), .ZN(n569) );
  OR2_X1 U652 ( .A1(n743), .A2(n569), .ZN(n572) );
  INV_X1 U653 ( .A(n570), .ZN(n571) );
  NAND2_X1 U654 ( .A1(n743), .A2(KEYINPUT44), .ZN(n574) );
  XNOR2_X1 U655 ( .A(n574), .B(KEYINPUT87), .ZN(n575) );
  INV_X1 U656 ( .A(n575), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n358), .A2(n578), .ZN(n651) );
  NOR2_X1 U658 ( .A1(n651), .A2(n584), .ZN(n580) );
  XNOR2_X1 U659 ( .A(n580), .B(n579), .ZN(n632) );
  OR2_X1 U660 ( .A1(n582), .A2(n358), .ZN(n583) );
  NOR2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT94), .ZN(n617) );
  NAND2_X1 U663 ( .A1(n353), .A2(n524), .ZN(n592) );
  INV_X1 U664 ( .A(n643), .ZN(n587) );
  NOR2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U667 ( .A(KEYINPUT102), .ZN(n593) );
  XNOR2_X1 U668 ( .A(n677), .B(KEYINPUT2), .ZN(n597) );
  INV_X1 U669 ( .A(n595), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n599) );
  INV_X1 U671 ( .A(KEYINPUT64), .ZN(n598) );
  XNOR2_X2 U672 ( .A(n599), .B(n598), .ZN(n697) );
  NAND2_X1 U673 ( .A1(n697), .A2(G472), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(n601), .ZN(n603) );
  NOR2_X2 U675 ( .A1(n603), .A2(n717), .ZN(n605) );
  INV_X1 U676 ( .A(KEYINPUT63), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n605), .B(n604), .ZN(G57) );
  XNOR2_X1 U678 ( .A(n606), .B(G119), .ZN(G21) );
  XNOR2_X1 U679 ( .A(n607), .B(G140), .ZN(G42) );
  NAND2_X1 U680 ( .A1(n697), .A2(G210), .ZN(n611) );
  XNOR2_X1 U681 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X2 U684 ( .A1(n612), .A2(n717), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U686 ( .A(G101), .B(n614), .Z(G3) );
  XOR2_X1 U687 ( .A(G104), .B(KEYINPUT107), .Z(n616) );
  NAND2_X1 U688 ( .A1(n628), .A2(n617), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(G6) );
  XOR2_X1 U690 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n619) );
  NAND2_X1 U691 ( .A1(n631), .A2(n617), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U693 ( .A(G107), .B(n620), .ZN(G9) );
  XNOR2_X1 U694 ( .A(G110), .B(n621), .ZN(G12) );
  XOR2_X1 U695 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U696 ( .A1(n631), .A2(n626), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(G30) );
  XNOR2_X1 U698 ( .A(n624), .B(G143), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT108), .B(n625), .ZN(G45) );
  NAND2_X1 U700 ( .A1(n626), .A2(n628), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(G146), .ZN(G48) );
  XOR2_X1 U702 ( .A(G113), .B(KEYINPUT109), .Z(n630) );
  NAND2_X1 U703 ( .A1(n632), .A2(n628), .ZN(n629) );
  XNOR2_X1 U704 ( .A(n630), .B(n629), .ZN(G15) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n633), .B(KEYINPUT110), .ZN(n634) );
  XNOR2_X1 U707 ( .A(G116), .B(n634), .ZN(G18) );
  XOR2_X1 U708 ( .A(G125), .B(KEYINPUT37), .Z(n635) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(G27) );
  XNOR2_X1 U710 ( .A(G134), .B(n637), .ZN(G36) );
  XNOR2_X1 U711 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n638), .B(KEYINPUT51), .ZN(n654) );
  INV_X1 U713 ( .A(n639), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(KEYINPUT50), .ZN(n650) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT49), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(KEYINPUT111), .B(n648), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U722 ( .A(n654), .B(n653), .Z(n655) );
  NOR2_X1 U723 ( .A1(n672), .A2(n655), .ZN(n666) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U728 ( .A1(n357), .A2(n664), .ZN(n665) );
  NOR2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U730 ( .A(n667), .B(KEYINPUT52), .ZN(n668) );
  XNOR2_X1 U731 ( .A(KEYINPUT114), .B(n668), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U733 ( .A(KEYINPUT115), .B(n671), .Z(n675) );
  NOR2_X1 U734 ( .A1(n357), .A2(n672), .ZN(n674) );
  NOR2_X1 U735 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U736 ( .A(n676), .B(KEYINPUT116), .ZN(n688) );
  BUF_X1 U737 ( .A(n677), .Z(n681) );
  INV_X1 U738 ( .A(n681), .ZN(n679) );
  NOR2_X1 U739 ( .A1(KEYINPUT2), .A2(KEYINPUT85), .ZN(n678) );
  NAND2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n683) );
  XNOR2_X1 U741 ( .A(KEYINPUT86), .B(KEYINPUT2), .ZN(n684) );
  OR2_X1 U742 ( .A1(n684), .A2(KEYINPUT85), .ZN(n680) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n686) );
  NAND2_X1 U745 ( .A1(n684), .A2(KEYINPUT85), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n689), .A2(n359), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n690), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U750 ( .A1(n711), .A2(G469), .ZN(n695) );
  XNOR2_X1 U751 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n693) );
  XNOR2_X1 U752 ( .A(n691), .B(KEYINPUT57), .ZN(n692) );
  XNOR2_X1 U753 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U754 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n717), .A2(n696), .ZN(G54) );
  NAND2_X1 U756 ( .A1(n697), .A2(G475), .ZN(n704) );
  XNOR2_X1 U757 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n698) );
  XNOR2_X1 U758 ( .A(n698), .B(KEYINPUT59), .ZN(n699) );
  XNOR2_X1 U759 ( .A(KEYINPUT90), .B(n699), .ZN(n702) );
  XNOR2_X1 U760 ( .A(n700), .B(KEYINPUT65), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n702), .B(n701), .ZN(n703) );
  INV_X1 U762 ( .A(n717), .ZN(n705) );
  XNOR2_X1 U763 ( .A(KEYINPUT60), .B(n707), .ZN(G60) );
  NAND2_X1 U764 ( .A1(n711), .A2(G478), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U766 ( .A1(n717), .A2(n710), .ZN(G63) );
  NAND2_X1 U767 ( .A1(n711), .A2(G217), .ZN(n715) );
  XOR2_X1 U768 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n712) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n359), .A2(G224), .ZN(n718) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n719), .A2(G898), .ZN(n720) );
  XOR2_X1 U773 ( .A(KEYINPUT122), .B(n720), .Z(n721) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n729) );
  XNOR2_X1 U775 ( .A(G101), .B(n723), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n724), .B(G110), .ZN(n726) );
  NOR2_X1 U777 ( .A1(G898), .A2(n733), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U779 ( .A(KEYINPUT123), .B(n727), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n729), .B(n728), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n730), .B(n731), .ZN(n736) );
  XOR2_X1 U782 ( .A(n736), .B(n732), .Z(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n735), .B(KEYINPUT124), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n736), .B(G227), .ZN(n737) );
  XNOR2_X1 U786 ( .A(n737), .B(KEYINPUT125), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n359), .A2(n739), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U790 ( .A(KEYINPUT126), .B(n742), .ZN(G72) );
  XOR2_X1 U791 ( .A(n743), .B(G122), .Z(G24) );
  XOR2_X1 U792 ( .A(n744), .B(G137), .Z(G39) );
  XOR2_X1 U793 ( .A(G131), .B(n745), .Z(G33) );
endmodule

