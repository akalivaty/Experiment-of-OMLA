//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT68), .B(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n463), .A3(G137), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G101), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n479), .B2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n466), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n463), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n479), .A2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n489), .A2(new_n491), .B1(new_n492), .B2(G136), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n488), .A2(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n464), .B2(new_n465), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n473), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n495), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n477), .C2(new_n478), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT71), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n481), .B(new_n483), .C1(new_n477), .C2(new_n478), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n466), .A2(new_n463), .A3(new_n510), .A4(G138), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n501), .A2(new_n506), .B1(new_n509), .B2(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n515), .B1(KEYINPUT6), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT72), .B(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(new_n516), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n515), .B(G651), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n514), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n514), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n525), .A2(G88), .B1(G651), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n524), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G50), .A3(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(G166));
  XNOR2_X1  g107(.A(KEYINPUT75), .B(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n537), .A2(new_n541), .B1(new_n513), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n530), .A2(G51), .A3(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(new_n525), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n530), .A2(G52), .A3(G543), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n516), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n525), .A2(G81), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n530), .A2(G43), .A3(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n514), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n525), .A2(G81), .B1(G651), .B2(new_n558), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n563), .A2(KEYINPUT76), .A3(new_n555), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(G860), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT77), .Z(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT78), .B(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n514), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n525), .A2(G91), .B1(G651), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  AND2_X1   g150(.A1(G53), .A2(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n530), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n575), .B1(new_n530), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n530), .A2(new_n576), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT9), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n577), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n585), .A2(KEYINPUT79), .A3(new_n574), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G299));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n544), .B2(new_n545), .ZN(new_n590));
  AND4_X1   g165(.A1(new_n589), .A2(new_n534), .A3(new_n543), .A4(new_n545), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(G286));
  NAND2_X1  g167(.A1(new_n529), .A2(new_n531), .ZN(G303));
  OAI21_X1  g168(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT81), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G87), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n530), .A2(G49), .A3(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  OAI21_X1  g173(.A(KEYINPUT73), .B1(new_n522), .B2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n599), .B1(new_n602), .B2(G651), .ZN(new_n603));
  AOI211_X1 g178(.A(KEYINPUT73), .B(new_n516), .C1(new_n600), .C2(new_n601), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G48), .A2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT82), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  INV_X1    g183(.A(new_n606), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n530), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n612));
  NAND2_X1  g187(.A1(G73), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G61), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n514), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n525), .A2(G86), .B1(G651), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n612), .B1(new_n611), .B2(new_n616), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(G305));
  NAND2_X1  g195(.A1(new_n525), .A2(G85), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G47), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n530), .A2(G543), .ZN(new_n624));
  OAI221_X1 g199(.A(new_n621), .B1(new_n516), .B2(new_n622), .C1(new_n623), .C2(new_n624), .ZN(G290));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(G301), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n530), .A2(G54), .A3(G543), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(new_n516), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n525), .A2(G92), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n627), .B1(new_n639), .B2(new_n626), .ZN(G284));
  XOR2_X1   g215(.A(G284), .B(KEYINPUT85), .Z(G321));
  MUX2_X1   g216(.A(G286), .B(G299), .S(new_n626), .Z(G297));
  MUX2_X1   g217(.A(G286), .B(G299), .S(new_n626), .Z(G280));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n639), .B1(new_n644), .B2(G860), .ZN(G148));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n646), .A3(new_n644), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n637), .A2(new_n638), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT86), .B1(new_n648), .B2(G559), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n626), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n562), .A2(new_n564), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n650), .A2(new_n651), .B1(new_n626), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n650), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g230(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT13), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n487), .A2(G123), .ZN(new_n661));
  INV_X1    g236(.A(G111), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n663));
  OAI21_X1  g238(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n484), .A2(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n663), .ZN(new_n666));
  AOI22_X1  g241(.A1(new_n665), .A2(new_n666), .B1(new_n492), .B2(G135), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(G2096), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n659), .A2(G2100), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(G2096), .ZN(new_n671));
  NAND4_X1  g246(.A1(new_n660), .A2(new_n669), .A3(new_n670), .A4(new_n671), .ZN(G156));
  XOR2_X1   g247(.A(G2451), .B(G2454), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT14), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2427), .B(G2438), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2430), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT15), .B(G2435), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n676), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(G2443), .B(G2446), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  AND3_X1   g261(.A1(new_n685), .A2(G14), .A3(new_n686), .ZN(G401));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT17), .ZN(new_n690));
  XOR2_X1   g265(.A(G2067), .B(G2678), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2084), .B(G2090), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n689), .B2(new_n692), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n690), .B2(new_n692), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n691), .A2(new_n693), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT18), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n694), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G2096), .B(G2100), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G227));
  XOR2_X1   g277(.A(G1971), .B(G1976), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT19), .ZN(new_n704));
  XOR2_X1   g279(.A(G1956), .B(G2474), .Z(new_n705));
  XOR2_X1   g280(.A(G1961), .B(G1966), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n704), .A2(new_n709), .A3(new_n707), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n712));
  AOI211_X1 g287(.A(new_n708), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT91), .Z(new_n715));
  XOR2_X1   g290(.A(G1981), .B(G1986), .Z(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n715), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G22), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1971), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT95), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n723), .A2(G23), .ZN(new_n728));
  INV_X1    g303(.A(G288), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n723), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT33), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1976), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G6), .B(G305), .S(G16), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT32), .B(G1981), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n733), .A2(new_n736), .A3(KEYINPUT34), .ZN(new_n737));
  MUX2_X1   g312(.A(G24), .B(G290), .S(G16), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT93), .B(G1986), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n742));
  NOR2_X1   g317(.A1(G25), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n487), .A2(G119), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n463), .A2(G107), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n745), .A2(new_n747), .B1(new_n492), .B2(G131), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT35), .B(G1991), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n751), .B(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n741), .A2(new_n742), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT34), .B1(new_n733), .B2(new_n736), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n737), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n737), .A2(new_n755), .A3(new_n759), .A4(new_n756), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n639), .A2(new_n723), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G4), .B2(new_n723), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n492), .A2(G139), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n770), .C1(new_n463), .C2(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G33), .B(new_n772), .S(G29), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2072), .ZN(new_n774));
  INV_X1    g349(.A(G29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n775), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT29), .B(G2090), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(G160), .A2(G29), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G34), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(new_n775), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n780), .A2(G2084), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(G2084), .B1(new_n780), .B2(new_n783), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT30), .B(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n786), .A2(new_n775), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n668), .B2(new_n775), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n784), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n775), .A2(G26), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT28), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n487), .A2(G128), .ZN(new_n794));
  INV_X1    g369(.A(G2104), .ZN(new_n795));
  INV_X1    g370(.A(G116), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n484), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G104), .A2(G2105), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT98), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n797), .A2(new_n799), .B1(new_n492), .B2(G140), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n793), .B1(new_n801), .B2(G29), .ZN(new_n802));
  INV_X1    g377(.A(G2067), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n774), .A2(new_n779), .A3(new_n791), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n775), .A2(G32), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n492), .A2(G141), .ZN(new_n807));
  NAND3_X1  g382(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT26), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G129), .B2(new_n487), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(new_n775), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT27), .B(G1996), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n775), .A2(G27), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G164), .B2(new_n775), .ZN(new_n817));
  INV_X1    g392(.A(G2078), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n723), .A2(G21), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G168), .B2(new_n723), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n723), .A2(G5), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G171), .B2(new_n723), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n822), .A2(G1966), .B1(new_n824), .B2(G1961), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n820), .B(new_n825), .C1(G1961), .C2(new_n824), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n767), .A2(new_n805), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(G1966), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT100), .Z(new_n829));
  AND2_X1   g404(.A1(new_n723), .A2(G19), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n652), .B2(G16), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT97), .B(G1341), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n723), .A2(G20), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT23), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n587), .B2(new_n723), .ZN(new_n838));
  INV_X1    g413(.A(G1956), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n765), .B2(new_n766), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n827), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n762), .A2(new_n763), .A3(new_n842), .ZN(G311));
  NAND3_X1  g418(.A1(new_n762), .A2(new_n763), .A3(new_n842), .ZN(G150));
  NAND2_X1  g419(.A1(new_n525), .A2(G93), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n530), .A2(G55), .A3(G543), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n516), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n562), .B2(new_n564), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n560), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n648), .A2(new_n644), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n851), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g438(.A(new_n812), .B(new_n801), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n502), .A2(new_n505), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n509), .B2(new_n511), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n864), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n772), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n487), .A2(G130), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT103), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n463), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n492), .B2(G142), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n492), .A2(KEYINPUT102), .A3(G142), .ZN(new_n875));
  OAI221_X1 g450(.A(new_n871), .B1(new_n872), .B2(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n749), .B(new_n657), .Z(new_n877));
  XOR2_X1   g452(.A(new_n876), .B(new_n877), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n869), .A2(KEYINPUT104), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n869), .B1(KEYINPUT104), .B2(new_n879), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n668), .B(G160), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(G162), .Z(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n869), .B2(new_n878), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n869), .B2(new_n878), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g464(.A1(G305), .A2(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(G290), .B(G303), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n729), .B1(new_n618), .B2(new_n619), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT42), .Z(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n647), .A2(new_n649), .ZN(new_n898));
  INV_X1    g473(.A(new_n853), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n647), .A2(new_n649), .A3(new_n853), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n582), .A2(new_n636), .A3(new_n586), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n636), .B1(new_n582), .B2(new_n586), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n900), .A2(new_n901), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n904), .A2(new_n905), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n900), .B2(new_n901), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n897), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n911), .ZN(new_n914));
  INV_X1    g489(.A(new_n901), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n853), .B1(new_n647), .B2(new_n649), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n900), .A2(new_n901), .A3(new_n909), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT105), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n896), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n896), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n851), .A2(new_n626), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(G331));
  NAND2_X1  g500(.A1(new_n546), .A2(G301), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(G286), .B2(G301), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n652), .A2(new_n851), .ZN(new_n928));
  INV_X1    g503(.A(new_n852), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(KEYINPUT106), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n850), .B2(new_n852), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n930), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n914), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n932), .ZN(new_n937));
  INV_X1    g512(.A(G286), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G171), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n939), .A3(new_n926), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n909), .A3(new_n933), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n941), .A3(new_n895), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n887), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n895), .B1(new_n936), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT108), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n940), .A2(new_n909), .A3(new_n933), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n911), .B1(new_n940), .B2(new_n933), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n895), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n936), .A2(new_n941), .A3(KEYINPUT107), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n942), .A2(new_n887), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n957), .B(KEYINPUT43), .C1(new_n943), .C2(new_n944), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n946), .A2(new_n956), .A3(KEYINPUT44), .A4(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n943), .A2(KEYINPUT43), .A3(new_n944), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n866), .B2(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(G160), .A2(G40), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n812), .B(G1996), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n801), .B(new_n803), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n749), .B(new_n752), .Z(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(G290), .B(G1986), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G8), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n509), .A2(new_n511), .ZN(new_n978));
  INV_X1    g553(.A(new_n865), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n471), .A2(new_n475), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(G288), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n983), .B(new_n988), .C1(new_n984), .C2(G288), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n987), .B(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n608), .B1(new_n530), .B2(new_n609), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT82), .B(new_n606), .C1(new_n519), .C2(new_n524), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n525), .A2(G86), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n615), .A2(G651), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(G1981), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n616), .B(new_n1000), .C1(new_n992), .C2(new_n993), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT115), .B(G1981), .C1(new_n994), .C2(new_n997), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n983), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n991), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT49), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(KEYINPUT116), .A3(new_n983), .A4(new_n1005), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n990), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n501), .A2(new_n506), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1021), .B2(new_n978), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n982), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT109), .ZN(new_n1025));
  NOR4_X1   g600(.A1(new_n866), .A2(KEYINPUT109), .A3(new_n965), .A4(G1384), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1023), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT110), .B(G1971), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(new_n978), .ZN(new_n1032));
  INV_X1    g607(.A(G1384), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g609(.A(new_n982), .B1(new_n980), .B2(new_n1031), .C1(new_n1034), .C2(KEYINPUT50), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1035), .A2(KEYINPUT118), .ZN(new_n1036));
  AOI21_X1  g611(.A(G2090), .B1(new_n1035), .B2(KEYINPUT118), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1020), .B1(new_n977), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n967), .B1(new_n980), .B2(new_n1031), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2090), .ZN(new_n1043));
  OAI221_X1 g618(.A(G8), .B1(new_n1030), .B2(new_n1043), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n966), .A2(new_n982), .ZN(new_n1046));
  NOR3_X1   g621(.A1(G164), .A2(new_n965), .A3(G1384), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n980), .A2(new_n1031), .ZN(new_n1049));
  INV_X1    g624(.A(G2084), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1041), .A2(new_n1049), .A3(new_n1050), .A4(new_n982), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n938), .A2(new_n1052), .A3(G8), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1012), .A2(new_n1039), .A3(new_n1044), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(KEYINPUT63), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1030), .B2(new_n1043), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1020), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(new_n1012), .A3(new_n1044), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1020), .A2(new_n1058), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1012), .A2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1012), .A2(new_n1039), .A3(new_n1044), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1048), .A2(G168), .A3(new_n1051), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  AND2_X1   g641(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(G8), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1052), .A2(G8), .A3(new_n546), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT62), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1068), .A2(new_n1075), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G2078), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1046), .A2(new_n1047), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(G1961), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n967), .B1(new_n1034), .B2(new_n965), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT109), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1082), .B(new_n818), .C1(new_n1084), .C2(new_n1026), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1080), .B(new_n1081), .C1(new_n1077), .C2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(G301), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1074), .A2(new_n1076), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1063), .B1(new_n1064), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G288), .A2(G1976), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT117), .B(new_n1001), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1001), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n983), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1061), .A2(new_n1089), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1996), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n980), .A2(KEYINPUT119), .A3(new_n982), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT119), .B1(new_n980), .B2(new_n982), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  AOI22_X1  g679(.A1(new_n1028), .A2(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n1105), .B2(new_n652), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1102), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n980), .A2(new_n982), .A3(KEYINPUT119), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1104), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1082), .B1(new_n1084), .B2(new_n1026), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(G1996), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n562), .A4(new_n564), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1042), .A2(new_n766), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n636), .A2(KEYINPUT60), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n803), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n636), .A2(KEYINPUT60), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1114), .A2(KEYINPUT60), .A3(new_n636), .A4(new_n1116), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1106), .A2(new_n1113), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1082), .B(new_n1122), .C1(new_n1084), .C2(new_n1026), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1034), .A2(KEYINPUT50), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n982), .B1(new_n980), .B2(new_n1031), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n839), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n574), .B(new_n1128), .C1(new_n578), .C2(new_n579), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n585), .B2(new_n574), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1123), .A2(new_n1132), .A3(new_n1126), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1126), .B2(new_n1123), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT61), .B1(new_n1138), .B2(KEYINPUT120), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(KEYINPUT121), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1123), .A2(new_n1132), .A3(new_n1142), .A4(new_n1126), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1141), .A2(new_n1143), .A3(KEYINPUT61), .A4(new_n1134), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1121), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1147));
  INV_X1    g722(.A(new_n636), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1134), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1136), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1145), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1081), .B1(new_n1085), .B2(new_n1077), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n467), .A2(new_n470), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n463), .B1(new_n1155), .B2(KEYINPUT124), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(KEYINPUT124), .B2(new_n1155), .ZN(new_n1157));
  INV_X1    g732(.A(new_n475), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1079), .A2(new_n981), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n966), .C1(new_n1084), .C2(new_n1026), .ZN(new_n1161));
  XOR2_X1   g736(.A(G301), .B(KEYINPUT54), .Z(new_n1162));
  NAND3_X1  g737(.A1(new_n1154), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1086), .B2(new_n1162), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1153), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1165), .A2(new_n1039), .A3(new_n1044), .A4(new_n1012), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1151), .A2(new_n1152), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n976), .B1(new_n1099), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n968), .A2(new_n1100), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT46), .ZN(new_n1170));
  INV_X1    g745(.A(new_n968), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n970), .A2(new_n812), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  OR3_X1    g749(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n974), .A2(new_n968), .B1(KEYINPUT48), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(KEYINPUT48), .B2(new_n1176), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n750), .A2(new_n752), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n971), .B2(new_n968), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n801), .A2(G2067), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1180), .A2(KEYINPUT125), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT125), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(new_n968), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1174), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT126), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1168), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g762(.A1(G227), .A2(new_n461), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  AND2_X1   g764(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  NOR4_X1   g766(.A1(G229), .A2(new_n1191), .A3(new_n1192), .A4(G401), .ZN(new_n1193));
  OAI211_X1 g767(.A(new_n888), .B(new_n1193), .C1(new_n961), .C2(new_n962), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


