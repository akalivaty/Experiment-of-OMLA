//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT69), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n453), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  INV_X1    g041(.A(G113), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n463), .B2(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(KEYINPUT70), .A3(new_n473), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n465), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n479), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g066(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n492));
  OAI221_X1 g067(.A(G2104), .B1(G112), .B2(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n498), .B(new_n500), .C1(new_n464), .C2(new_n463), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n489), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n489), .A2(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n477), .B2(new_n478), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n501), .B(new_n503), .C1(new_n505), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(G126), .A2(G2105), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n479), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g090(.A(KEYINPUT72), .B(new_n512), .C1(new_n463), .C2(new_n464), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(KEYINPUT6), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(KEYINPUT74), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n521), .A2(new_n522), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n528), .A2(KEYINPUT6), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(G88), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n532), .A2(G50), .A3(G543), .A4(new_n534), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n537), .B1(new_n535), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n526), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G166));
  NAND2_X1  g116(.A1(new_n532), .A2(new_n534), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n523), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n529), .A2(new_n531), .B1(KEYINPUT6), .B2(new_n528), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G51), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n550));
  AND2_X1   g125(.A1(G63), .A2(G651), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n549), .A2(new_n550), .B1(new_n533), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n544), .A2(new_n547), .A3(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  NAND2_X1  g129(.A1(new_n543), .A2(G90), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT76), .B(G52), .Z(new_n556));
  NAND2_X1  g131(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n533), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n528), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n523), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  XOR2_X1   g140(.A(KEYINPUT77), .B(G43), .Z(new_n566));
  NAND3_X1  g141(.A1(new_n545), .A2(G543), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n545), .A2(G81), .A3(new_n533), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT78), .Z(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g147(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n573));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(KEYINPUT80), .B2(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n546), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n545), .A2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n577), .B(new_n578), .C1(new_n583), .C2(new_n580), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n533), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n528), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n545), .A2(G91), .A3(new_n533), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n582), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n540), .A2(KEYINPUT81), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n590), .B(new_n526), .C1(new_n538), .C2(new_n539), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(G303));
  NAND4_X1  g167(.A1(new_n532), .A2(G87), .A3(new_n533), .A4(new_n534), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT82), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n545), .A2(new_n595), .A3(G87), .A4(new_n533), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n532), .A2(G49), .A3(G543), .A4(new_n534), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n597), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G288));
  NAND3_X1  g181(.A1(new_n545), .A2(G48), .A3(G543), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n545), .A2(G86), .A3(new_n533), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n521), .B2(new_n522), .ZN(new_n610));
  AND2_X1   g185(.A1(G73), .A2(G543), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(new_n543), .A2(G85), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n546), .A2(G47), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n533), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n614), .B(new_n615), .C1(new_n528), .C2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n523), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n546), .A2(G54), .B1(new_n621), .B2(G651), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n532), .A2(G92), .A3(new_n533), .A4(new_n534), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT10), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n624), .A2(KEYINPUT84), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(KEYINPUT84), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n623), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n618), .B1(new_n631), .B2(G868), .ZN(G284));
  OAI21_X1  g207(.A(new_n618), .B1(new_n631), .B2(G868), .ZN(G321));
  NAND2_X1  g208(.A1(G286), .A2(G868), .ZN(new_n634));
  AND4_X1   g209(.A1(new_n582), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G868), .ZN(G297));
  OAI21_X1  g211(.A(new_n634), .B1(new_n635), .B2(G868), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n631), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n631), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n479), .A2(new_n470), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT85), .B(KEYINPUT13), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n484), .A2(G135), .ZN(new_n649));
  INV_X1    g224(.A(G123), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n489), .A2(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  OAI221_X1 g227(.A(new_n649), .B1(new_n650), .B2(new_n487), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(G2096), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(G2096), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n648), .A2(new_n656), .A3(new_n657), .ZN(G156));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT87), .B(G2438), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR3_X1    g240(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(KEYINPUT14), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XOR2_X1   g245(.A(G1341), .B(G1348), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n672), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT18), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n681), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n682), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n680), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n684), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G2096), .B(G2100), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1956), .B(G2474), .Z(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n705), .B(new_n704), .S(new_n697), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(G229));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G168), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1966), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT100), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(G1966), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT102), .Z(new_n721));
  NOR2_X1   g296(.A1(G5), .A2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT103), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G301), .B2(new_n715), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT101), .B1(new_n655), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT30), .B(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n730), .A2(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  OR4_X1    g309(.A1(new_n719), .A2(new_n721), .A3(new_n726), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n715), .A2(G4), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n631), .B2(new_n715), .ZN(new_n739));
  INV_X1    g314(.A(G1348), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n484), .A2(G139), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n489), .A2(G103), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(new_n489), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT99), .ZN(new_n750));
  MUX2_X1   g325(.A(G33), .B(new_n750), .S(G29), .Z(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G2072), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n727), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n727), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT29), .Z(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(new_n725), .B2(new_n724), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n715), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT23), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n635), .B2(new_n715), .ZN(new_n760));
  INV_X1    g335(.A(G1956), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n752), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n715), .A2(G19), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT98), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n569), .B2(new_n715), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1341), .ZN(new_n767));
  NAND2_X1  g342(.A1(G164), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G27), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n727), .A2(G32), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n773));
  INV_X1    g348(.A(new_n487), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT26), .Z(new_n777));
  NAND3_X1  g352(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(new_n727), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n769), .A2(new_n770), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n484), .A2(G140), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n489), .ZN(new_n786));
  INV_X1    g361(.A(G128), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n786), .C1(new_n787), .C2(new_n487), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n727), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n771), .A2(new_n782), .A3(new_n783), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G34), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(KEYINPUT24), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(KEYINPUT24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n727), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G160), .B2(new_n727), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G2084), .Z(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n755), .B2(new_n756), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n763), .A2(new_n767), .A3(new_n795), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n736), .A2(new_n737), .A3(new_n741), .A4(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G25), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n805), .A2(KEYINPUT91), .A3(G29), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT91), .B1(new_n805), .B2(G29), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT93), .B1(G95), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(KEYINPUT93), .A2(G95), .A3(G2105), .ZN(new_n810));
  OAI221_X1 g385(.A(G2104), .B1(G107), .B2(new_n489), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT94), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n484), .A2(G131), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n774), .A2(G119), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n806), .B(new_n807), .C1(new_n816), .C2(new_n727), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  MUX2_X1   g394(.A(G24), .B(G290), .S(G16), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G305), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G16), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G6), .B2(G16), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT32), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(KEYINPUT32), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G1981), .ZN(new_n829));
  INV_X1    g404(.A(G1981), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G16), .A2(G22), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G166), .B2(G16), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT96), .B(G1971), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n601), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n597), .A2(KEYINPUT95), .A3(new_n600), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  MUX2_X1   g415(.A(G23), .B(new_n840), .S(G16), .Z(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT33), .B(G1976), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n843), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n832), .A2(new_n836), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n822), .B1(new_n846), .B2(KEYINPUT34), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT97), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n822), .B(new_n849), .C1(new_n846), .C2(KEYINPUT34), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT36), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n804), .B1(new_n854), .B2(new_n856), .ZN(G311));
  INV_X1    g432(.A(new_n804), .ZN(new_n858));
  INV_X1    g433(.A(new_n856), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n855), .B1(new_n851), .B2(new_n852), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(G150));
  NAND2_X1  g436(.A1(new_n631), .A2(G559), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT38), .Z(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  INV_X1    g439(.A(G67), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n523), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G651), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n545), .A2(G93), .A3(new_n533), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n545), .A2(G55), .A3(G543), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n863), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n876));
  AOI21_X1  g451(.A(G860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(G860), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT37), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G145));
  NAND2_X1  g456(.A1(new_n484), .A2(G142), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  INV_X1    g459(.A(G118), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(G2105), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n884), .B2(new_n883), .ZN(new_n887));
  INV_X1    g462(.A(G130), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n882), .B(new_n887), .C1(new_n888), .C2(new_n487), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT106), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n645), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n816), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n518), .B(new_n788), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n778), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n748), .B2(new_n746), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n750), .B2(new_n895), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n655), .B(new_n495), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n482), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n897), .B(new_n892), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n900), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(G395));
  XOR2_X1   g484(.A(new_n640), .B(new_n874), .Z(new_n910));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n631), .B2(G299), .ZN(new_n911));
  INV_X1    g486(.A(new_n630), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n628), .B1(new_n627), .B2(new_n629), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n622), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n635), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n631), .A2(G299), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n911), .A2(new_n916), .A3(new_n921), .A4(new_n917), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n923), .B2(new_n910), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n840), .B(new_n540), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(G305), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI221_X1 g507(.A(new_n919), .B1(new_n930), .B2(new_n931), .C1(new_n923), .C2(new_n910), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n925), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n925), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n867), .A2(new_n869), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n937), .A2(new_n868), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(G868), .B2(new_n938), .ZN(G295));
  OAI21_X1  g514(.A(new_n936), .B1(G868), .B2(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  OAI21_X1  g517(.A(G171), .B1(new_n872), .B2(new_n873), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n569), .A2(new_n868), .A3(new_n937), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n870), .A2(new_n871), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(G301), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n943), .A2(new_n946), .A3(G168), .ZN(new_n947));
  AOI21_X1  g522(.A(G168), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n918), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n920), .A2(new_n952), .A3(new_n922), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n918), .B(KEYINPUT109), .C1(new_n947), .C2(new_n948), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n951), .A2(new_n953), .A3(new_n928), .A4(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(new_n903), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n929), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n942), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n929), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n903), .A3(new_n955), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n941), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n941), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n956), .A2(new_n942), .A3(new_n958), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n965), .A2(KEYINPUT110), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT110), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G397));
  AOI21_X1  g544(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n467), .A2(new_n468), .ZN(new_n971));
  OAI21_X1  g546(.A(G2105), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n470), .A2(G101), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT111), .B(G40), .Z(new_n974));
  NAND4_X1  g549(.A1(new_n481), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n471), .A2(new_n977), .A3(new_n481), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n511), .B2(new_n517), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(G1996), .A3(new_n778), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT113), .Z(new_n984));
  XNOR2_X1  g559(.A(new_n788), .B(new_n793), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(G1996), .B2(new_n778), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n816), .B(new_n818), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT48), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n818), .A2(new_n984), .A3(new_n816), .A4(new_n987), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n788), .A2(G2067), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n982), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n982), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT46), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n985), .A2(new_n779), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n982), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n994), .A2(new_n997), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n979), .B2(new_n981), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n823), .A2(new_n830), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1010), .A2(KEYINPUT49), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT49), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n838), .A2(G1976), .A3(new_n839), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1009), .A2(new_n1014), .B1(new_n1016), .B2(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n979), .A2(new_n981), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1015), .A2(G8), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n602), .A2(new_n1021), .A3(new_n604), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1009), .A2(new_n1015), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(KEYINPUT116), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1017), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G1384), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT72), .B1(new_n479), .B2(new_n512), .ZN(new_n1031));
  INV_X1    g606(.A(new_n516), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1033), .B2(new_n510), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1033), .B2(new_n510), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1034), .A2(KEYINPUT114), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n979), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1971), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n976), .A2(new_n978), .B1(new_n981), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n981), .B2(new_n1042), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1036), .A2(new_n1045), .A3(KEYINPUT50), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n756), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1008), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n589), .A2(G8), .A3(new_n591), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n589), .A2(KEYINPUT55), .A3(G8), .A4(new_n591), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT118), .B1(new_n1028), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(new_n1008), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1020), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1026), .A2(KEYINPUT116), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1058), .A2(new_n1059), .A3(new_n1062), .A4(new_n1017), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT117), .B(G2084), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1966), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1034), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n980), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1008), .B(G286), .C1(new_n1066), .C2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1064), .A2(KEYINPUT63), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1055), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n981), .A2(new_n1042), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1036), .A2(KEYINPUT50), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n979), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1077), .A2(new_n756), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1056), .B1(new_n1078), .B2(new_n1008), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(new_n1062), .A3(new_n1017), .A4(new_n1064), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1070), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1073), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1072), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1044), .A2(new_n979), .A3(new_n1074), .A4(new_n1046), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1043), .A2(KEYINPUT120), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n725), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(G2078), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n980), .A2(new_n1068), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1037), .A2(new_n1038), .A3(new_n770), .A4(new_n979), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1091), .B1(new_n1092), .B2(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1080), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n1008), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G168), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1066), .A2(new_n1069), .A3(G286), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1066), .A2(new_n1069), .A3(G168), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT51), .B1(new_n1105), .B2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(KEYINPUT62), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1096), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1028), .A2(new_n1064), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n1021), .A3(new_n605), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1010), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1009), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1083), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1119));
  AND3_X1   g694(.A1(G160), .A2(G40), .A3(new_n1090), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1119), .A2(new_n1120), .B1(new_n1092), .B2(new_n1089), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1088), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1122), .B2(G171), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(G171), .B2(new_n1094), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1080), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1107), .A4(new_n1104), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1086), .A2(new_n740), .A3(new_n1087), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n979), .A2(new_n793), .A3(new_n981), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n914), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n631), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n914), .A3(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1133), .B2(KEYINPUT60), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n569), .B1(KEYINPUT121), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1019), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1037), .A2(new_n1038), .A3(new_n998), .A4(new_n979), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1142), .B(new_n1136), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1076), .A2(new_n761), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1148));
  XNOR2_X1  g723(.A(G299), .B(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT56), .B(G2072), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1037), .A2(new_n1038), .A3(new_n979), .A4(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1149), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1152), .A2(new_n1153), .A3(KEYINPUT61), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n635), .B(new_n1148), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1151), .ZN(new_n1157));
  AOI21_X1  g732(.A(G1956), .B1(new_n1043), .B2(new_n1075), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1155), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1146), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1146), .B(new_n1164), .C1(new_n1154), .C2(new_n1161), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1134), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1131), .A2(new_n1152), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n1153), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1126), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1122), .B2(G171), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1088), .A2(new_n1121), .A3(KEYINPUT123), .A4(G301), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n1095), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1118), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT124), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n1176), .A3(new_n1118), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1117), .B1(new_n1169), .B2(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n982), .B1(new_n991), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n990), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1007), .B1(new_n1179), .B2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g758(.A1(G227), .A2(new_n461), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1185), .B1(new_n677), .B2(new_n678), .ZN(new_n1186));
  OR2_X1    g760(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1187));
  AND2_X1   g761(.A1(new_n713), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1189));
  OAI211_X1 g763(.A(new_n1188), .B(new_n1189), .C1(new_n904), .C2(new_n906), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n959), .A2(new_n963), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1190), .A2(new_n1191), .ZN(G308));
  OR2_X1    g766(.A1(new_n1190), .A2(new_n1191), .ZN(G225));
endmodule


