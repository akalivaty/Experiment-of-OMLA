//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n866, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  XNOR2_X1  g000(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT69), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(G120gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n203), .A2(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n203), .B2(G120gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G127gat), .ZN(new_n214));
  INV_X1    g013(.A(G127gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G134gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G113gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n208), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT67), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  INV_X1    g029(.A(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR3_X1   g037(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n236), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G155gat), .ZN(new_n241));
  INV_X1    g040(.A(G162gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n233), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n236), .ZN(new_n244));
  AND2_X1   g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT76), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n248), .A3(new_n234), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n220), .A2(new_n228), .A3(new_n240), .A4(new_n250), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n202), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n250), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n260), .A3(new_n229), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n240), .A2(new_n250), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n228), .A4(new_n220), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n261), .A2(new_n263), .A3(new_n265), .A4(new_n255), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n257), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n202), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n220), .A2(new_n228), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n264), .A3(new_n262), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n253), .A2(KEYINPUT4), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n261), .A2(new_n255), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT80), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(KEYINPUT6), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n275), .B2(new_n282), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n266), .A2(new_n257), .B1(new_n272), .B2(new_n273), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT28), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n300), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302));
  INV_X1    g101(.A(G169gat), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n298), .A2(new_n299), .A3(new_n301), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n296), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n321), .A3(new_n299), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n316), .A2(KEYINPUT64), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n316), .A2(KEYINPUT64), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n315), .A3(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n324), .A2(new_n325), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n269), .B1(new_n312), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n295), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n294), .B1(new_n290), .B2(new_n291), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n307), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT66), .B1(new_n306), .B2(new_n307), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n326), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n317), .A2(new_n313), .A3(new_n314), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n325), .B1(new_n339), .B2(new_n322), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n341), .A3(new_n229), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n331), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT34), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT34), .ZN(new_n346));
  INV_X1    g145(.A(new_n344), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n346), .B(new_n347), .C1(new_n331), .C2(new_n342), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT71), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n337), .A2(new_n229), .A3(new_n341), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n229), .B1(new_n337), .B2(new_n341), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n346), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(KEYINPUT34), .A3(new_n344), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n331), .A2(new_n347), .A3(new_n342), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT33), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n364), .B2(KEYINPUT33), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n360), .A2(new_n364), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n356), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n353), .A2(new_n355), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n363), .B1(new_n357), .B2(new_n359), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n357), .A2(new_n365), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n368), .B(KEYINPUT71), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT36), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT36), .B1(new_n367), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  INV_X1    g175(.A(G218gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(G197gat), .A2(G204gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n375), .B(new_n378), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n382), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n384), .B(new_n385), .C1(new_n380), .C2(new_n379), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT72), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n312), .A2(new_n330), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n337), .A2(new_n341), .B1(new_n392), .B2(new_n389), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n387), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n312), .A2(new_n330), .B1(KEYINPUT29), .B2(new_n390), .ZN(new_n395));
  INV_X1    g194(.A(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n337), .A2(new_n341), .A3(new_n389), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT74), .ZN(new_n400));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT30), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n394), .A2(new_n398), .A3(new_n405), .A4(new_n402), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT73), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n391), .A2(new_n393), .A3(new_n387), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n396), .B1(new_n395), .B2(new_n397), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n398), .A3(KEYINPUT73), .ZN(new_n412));
  INV_X1    g211(.A(new_n402), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n288), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n383), .B2(new_n386), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n251), .B1(new_n417), .B2(KEYINPUT3), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n260), .A2(new_n392), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n387), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n422), .B(new_n418), .C1(new_n419), .C2(new_n416), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(KEYINPUT83), .B(G22gat), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429));
  INV_X1    g228(.A(new_n427), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(new_n430), .A3(new_n425), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT31), .ZN(new_n434));
  INV_X1    g233(.A(G50gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT81), .Z(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n424), .B2(new_n425), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(G22gat), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n428), .B(new_n441), .C1(new_n442), .C2(new_n426), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n415), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n275), .A2(KEYINPUT85), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n267), .A2(new_n274), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n281), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n283), .B1(new_n449), .B2(new_n285), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n411), .A2(KEYINPUT37), .A3(new_n412), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n394), .A2(new_n398), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n454), .A2(new_n413), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT37), .B1(new_n409), .B2(new_n410), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(new_n451), .A3(new_n413), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n403), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n450), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n443), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n407), .A2(new_n414), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n267), .A2(new_n274), .A3(new_n447), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n447), .B1(new_n267), .B2(new_n274), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n282), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n270), .A2(new_n271), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n255), .B1(new_n466), .B2(new_n261), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT39), .B1(new_n254), .B2(new_n256), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n281), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  INV_X1    g272(.A(new_n471), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n281), .B1(new_n467), .B2(new_n468), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n374), .B(new_n445), .C1(new_n460), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n367), .A2(new_n371), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT35), .B1(new_n481), .B2(new_n415), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n371), .A2(new_n367), .B1(new_n440), .B2(new_n443), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n450), .A4(new_n462), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT88), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  OR2_X1    g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(G43gat), .A2(G50gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(G29gat), .A2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(KEYINPUT90), .A2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(KEYINPUT90), .A2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G29gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n493), .A2(new_n492), .A3(new_n494), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n496), .A2(new_n499), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n497), .B(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n500), .B2(new_n501), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n495), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  INV_X1    g311(.A(G1gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT16), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(G1gat), .B1(new_n511), .B2(KEYINPUT91), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n516), .A2(new_n517), .A3(G8gat), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n511), .A2(KEYINPUT91), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n521), .B2(new_n515), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n510), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n509), .A3(KEYINPUT17), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n519), .A3(new_n515), .ZN(new_n525));
  OAI21_X1  g324(.A(G8gat), .B1(new_n516), .B2(new_n517), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT17), .B1(new_n505), .B2(new_n509), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n491), .B(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT12), .ZN(new_n537));
  INV_X1    g336(.A(new_n528), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n518), .A2(new_n522), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(new_n524), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n491), .A4(new_n523), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n509), .A4(new_n505), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n491), .B(KEYINPUT13), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n531), .A2(new_n537), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n529), .A2(new_n530), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(KEYINPUT92), .A3(new_n541), .A4(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n541), .ZN(new_n552));
  INV_X1    g351(.A(new_n537), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n488), .A2(new_n490), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT93), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n488), .A2(new_n558), .A3(new_n490), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  XOR2_X1   g360(.A(G57gat), .B(G64gat), .Z(new_n562));
  OR2_X1    g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n564), .B(new_n563), .C1(new_n569), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n539), .B1(new_n561), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G183gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT94), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n573), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n561), .ZN(new_n579));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n376), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n590), .A2(new_n591), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n593), .A3(new_n587), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n599), .A2(new_n510), .B1(KEYINPUT41), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT97), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n524), .A2(new_n598), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n601), .B(new_n603), .C1(new_n604), .C2(new_n528), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT95), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n600), .A2(KEYINPUT41), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n601), .B1(new_n528), .B2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(new_n603), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(KEYINPUT98), .A3(new_n612), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n609), .B(KEYINPUT96), .Z(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n613), .B2(new_n605), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n583), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G176gat), .ZN(new_n625));
  INV_X1    g424(.A(G204gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT102), .Z(new_n630));
  NOR2_X1   g429(.A1(new_n592), .A2(new_n594), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n593), .B1(new_n596), .B2(new_n587), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n571), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n595), .A2(new_n597), .A3(new_n570), .A4(new_n568), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n571), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n630), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT103), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n628), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n636), .A2(new_n638), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n636), .B2(new_n638), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n629), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n645), .A3(new_n627), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n647), .A2(KEYINPUT104), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT104), .B1(new_n647), .B2(new_n652), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n623), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n560), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n659), .B(new_n656), .C1(new_n557), .C2(new_n559), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n289), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g461(.A1(new_n407), .A2(new_n414), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  OAI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n658), .C2(new_n660), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n479), .A2(new_n489), .A3(new_n486), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n489), .B1(new_n479), .B2(new_n486), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n558), .B1(new_n670), .B2(new_n555), .ZN(new_n671));
  INV_X1    g470(.A(new_n559), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n657), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n659), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n560), .A2(KEYINPUT105), .A3(new_n657), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n663), .A4(new_n664), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n663), .B1(new_n658), .B2(new_n660), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G8gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n667), .A2(new_n677), .A3(new_n679), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n676), .A2(new_n681), .A3(new_n480), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n372), .B2(new_n373), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n480), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT36), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n674), .B2(new_n675), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n682), .B1(new_n681), .B2(new_n690), .ZN(G1326gat));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT107), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n676), .B2(new_n444), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n444), .B(new_n693), .C1(new_n658), .C2(new_n660), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(G1327gat));
  NAND3_X1  g496(.A1(new_n655), .A2(new_n583), .A3(new_n622), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n560), .A2(new_n507), .A3(new_n289), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n488), .A2(KEYINPUT44), .A3(new_n490), .A4(new_n622), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  INV_X1    g504(.A(new_n477), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n444), .B1(new_n706), .B2(new_n663), .ZN(new_n707));
  INV_X1    g506(.A(new_n285), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n465), .A2(new_n708), .B1(KEYINPUT6), .B2(new_n287), .ZN(new_n709));
  INV_X1    g508(.A(new_n459), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n452), .A2(new_n455), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n709), .B(new_n710), .C1(new_n451), .C2(new_n711), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n707), .A2(new_n712), .B1(new_n444), .B2(new_n415), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n689), .A2(new_n713), .B1(new_n482), .B2(new_n485), .ZN(new_n714));
  INV_X1    g513(.A(new_n622), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n705), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n704), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n655), .ZN(new_n718));
  INV_X1    g517(.A(new_n583), .ZN(new_n719));
  INV_X1    g518(.A(new_n555), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n717), .A2(new_n289), .A3(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n702), .B(new_n703), .C1(new_n507), .C2(new_n722), .ZN(G1328gat));
  INV_X1    g522(.A(new_n502), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n560), .A2(new_n663), .A3(new_n724), .A4(new_n699), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n717), .A2(new_n663), .A3(new_n721), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n726), .A2(new_n727), .B1(new_n502), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT108), .B1(new_n726), .B2(new_n727), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n725), .A2(new_n731), .A3(KEYINPUT46), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734));
  INV_X1    g533(.A(new_n480), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n560), .A2(new_n699), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738));
  INV_X1    g537(.A(new_n689), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n704), .A2(new_n716), .A3(new_n739), .A4(new_n721), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n738), .B1(new_n737), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n734), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(G1330gat));
  NAND3_X1  g548(.A1(new_n717), .A2(new_n444), .A3(new_n721), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G50gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n560), .A2(new_n435), .A3(new_n444), .A4(new_n699), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1331gat));
  INV_X1    g554(.A(new_n714), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n720), .A3(new_n623), .A4(new_n718), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n289), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g560(.A(new_n757), .B(KEYINPUT110), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n462), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n762), .A2(G71gat), .A3(new_n735), .ZN(new_n769));
  INV_X1    g568(.A(G71gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n759), .B2(new_n739), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G71gat), .B1(new_n762), .B2(new_n689), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n759), .A2(new_n770), .A3(new_n480), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(KEYINPUT50), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n444), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n719), .A2(new_n555), .A3(new_n655), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n717), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n289), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n714), .A2(new_n715), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n719), .A2(new_n555), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n783), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(KEYINPUT111), .A3(new_n785), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n718), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n289), .A2(new_n585), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n781), .A2(new_n585), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n717), .A2(new_n663), .A3(new_n779), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n462), .A2(G92gat), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n794), .B(new_n796), .C1(new_n791), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n786), .A2(KEYINPUT112), .A3(new_n788), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n782), .B2(new_n783), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n655), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n796), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n799), .B1(new_n805), .B2(new_n794), .ZN(G1337gat));
  NAND2_X1  g605(.A1(new_n780), .A2(new_n739), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n655), .A2(new_n735), .A3(G99gat), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT113), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n790), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1338gat));
  NOR2_X1   g611(.A1(new_n461), .A2(G106gat), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n789), .A2(new_n718), .A3(new_n790), .A4(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n717), .A2(new_n444), .A3(new_n779), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G106gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n803), .A3(new_n813), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n817), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n627), .B1(new_n640), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n636), .A2(new_n638), .ZN(new_n825));
  INV_X1    g624(.A(new_n630), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n822), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n651), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT55), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT103), .B1(new_n825), .B2(new_n826), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT103), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n832), .B(new_n630), .C1(new_n636), .C2(new_n638), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n822), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n829), .A2(new_n834), .A3(KEYINPUT55), .A4(new_n628), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n829), .A2(new_n628), .A3(new_n834), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n646), .A2(new_n628), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n551), .A2(new_n554), .B1(new_n651), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n491), .B1(new_n540), .B2(new_n523), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n543), .A2(new_n544), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n536), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n551), .B(new_n846), .C1(new_n653), .C2(new_n654), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n622), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n652), .B1(new_n617), .B2(new_n620), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n839), .B2(new_n838), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n551), .A2(new_n846), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n551), .A2(KEYINPUT115), .A3(new_n846), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n837), .A2(new_n850), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n583), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n623), .A2(new_n720), .A3(new_n655), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n288), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n663), .A3(new_n481), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n555), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n204), .B2(new_n206), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n203), .B2(new_n861), .ZN(G1340gat));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n718), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n719), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(G127gat), .ZN(G1342gat));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n860), .B(new_n622), .C1(new_n868), .C2(new_n213), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n213), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(G1343gat));
  XNOR2_X1  g670(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n739), .A2(new_n288), .A3(new_n663), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n829), .A2(new_n834), .A3(new_n876), .A4(new_n628), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n839), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n837), .A2(new_n878), .A3(new_n842), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n622), .B1(new_n879), .B2(new_n847), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n583), .B1(new_n880), .B2(new_n855), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n874), .B(new_n461), .C1(new_n881), .C2(new_n857), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n461), .B1(new_n856), .B2(new_n857), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n882), .A2(new_n883), .B1(KEYINPUT57), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n857), .ZN(new_n886));
  AND4_X1   g685(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT57), .A4(new_n444), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n555), .B(new_n873), .C1(new_n885), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n689), .A2(new_n462), .A3(new_n444), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n858), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n555), .A2(new_n230), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT119), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n890), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n872), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n872), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n899), .B(new_n896), .C1(new_n888), .C2(G141gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(G1344gat));
  AND2_X1   g700(.A1(new_n890), .A2(new_n893), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n231), .A3(new_n718), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n873), .B1(new_n885), .B2(new_n887), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n655), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n884), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n886), .A2(new_n874), .A3(new_n444), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n718), .A3(new_n873), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n906), .B1(new_n913), .B2(G148gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n903), .B1(new_n908), .B2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n904), .B2(new_n583), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n902), .A2(new_n241), .A3(new_n719), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1346gat));
  OAI21_X1  g717(.A(G162gat), .B1(new_n904), .B2(new_n715), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n242), .A3(new_n622), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n856), .A2(new_n857), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n663), .A2(new_n288), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n481), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n303), .A3(new_n720), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(KEYINPUT121), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n555), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(new_n303), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n304), .A3(new_n718), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n925), .B2(new_n655), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1349gat));
  AND2_X1   g731(.A1(new_n922), .A2(new_n924), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n290), .A3(new_n719), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n933), .A2(KEYINPUT122), .A3(new_n290), .A4(new_n719), .ZN(new_n937));
  OAI21_X1  g736(.A(G183gat), .B1(new_n925), .B2(new_n583), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n940));
  NAND2_X1  g739(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT124), .Z(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n939), .B(new_n942), .C1(KEYINPUT123), .C2(KEYINPUT60), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n925), .B2(new_n715), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n927), .A2(new_n291), .A3(new_n622), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1351gat));
  NAND3_X1  g749(.A1(new_n689), .A2(new_n288), .A3(new_n663), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n910), .A2(new_n911), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n555), .A2(G197gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n909), .A2(new_n720), .A3(new_n951), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n953), .A2(new_n954), .B1(G197gat), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT125), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n909), .A2(new_n951), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n626), .A3(new_n718), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT126), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n958), .A2(new_n962), .A3(new_n626), .A4(new_n718), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT127), .Z(new_n964));
  NAND3_X1  g763(.A1(new_n912), .A2(new_n718), .A3(new_n952), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n376), .A3(new_n719), .ZN(new_n968));
  OAI21_X1  g767(.A(G211gat), .B1(new_n953), .B2(new_n583), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  NOR3_X1   g772(.A1(new_n953), .A2(new_n377), .A3(new_n715), .ZN(new_n974));
  AOI21_X1  g773(.A(G218gat), .B1(new_n958), .B2(new_n622), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(G1355gat));
endmodule


