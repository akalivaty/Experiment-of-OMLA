

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586;

  XNOR2_X1 U320 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U321 ( .A(n448), .B(KEYINPUT125), .ZN(n449) );
  XNOR2_X1 U322 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n445) );
  XNOR2_X1 U323 ( .A(n446), .B(n445), .ZN(n570) );
  XNOR2_X1 U324 ( .A(n399), .B(n398), .ZN(n404) );
  XNOR2_X1 U325 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U326 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U327 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U328 ( .A(G43GAT), .B(G134GAT), .Z(n356) );
  XNOR2_X1 U329 ( .A(G99GAT), .B(G71GAT), .ZN(n288) );
  XNOR2_X1 U330 ( .A(n288), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U331 ( .A(n356), .B(n402), .ZN(n289) );
  XOR2_X1 U332 ( .A(G15GAT), .B(G127GAT), .Z(n417) );
  XNOR2_X1 U333 ( .A(n289), .B(n417), .ZN(n290) );
  XOR2_X1 U334 ( .A(G113GAT), .B(KEYINPUT0), .Z(n331) );
  XOR2_X1 U335 ( .A(n290), .B(n331), .Z(n292) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U338 ( .A(KEYINPUT82), .B(KEYINPUT79), .Z(n294) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n296), .B(n295), .Z(n303) );
  XOR2_X1 U342 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n298) );
  XNOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(n299), .B(G183GAT), .Z(n301) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(G176GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n434) );
  XNOR2_X1 U348 ( .A(n434), .B(KEYINPUT80), .ZN(n302) );
  XOR2_X1 U349 ( .A(n303), .B(n302), .Z(n498) );
  INV_X1 U350 ( .A(n498), .ZN(n533) );
  XOR2_X1 U351 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT22), .B(KEYINPUT84), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U354 ( .A(G204GAT), .B(KEYINPUT85), .Z(n307) );
  XOR2_X1 U355 ( .A(G50GAT), .B(G162GAT), .Z(n347) );
  XOR2_X1 U356 ( .A(G22GAT), .B(G155GAT), .Z(n409) );
  XNOR2_X1 U357 ( .A(n347), .B(n409), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U359 ( .A(n309), .B(n308), .Z(n311) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n314) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n313) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n332) );
  XOR2_X1 U365 ( .A(n314), .B(n332), .Z(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n316) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G211GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n318) );
  XOR2_X1 U369 ( .A(G218GAT), .B(KEYINPUT86), .Z(n317) );
  XOR2_X1 U370 ( .A(n318), .B(n317), .Z(n442) );
  INV_X1 U371 ( .A(n442), .ZN(n320) );
  XNOR2_X1 U372 ( .A(G106GAT), .B(G78GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n319), .B(G148GAT), .ZN(n393) );
  XOR2_X1 U374 ( .A(n320), .B(n393), .Z(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n466) );
  XOR2_X1 U376 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n324) );
  XNOR2_X1 U377 ( .A(KEYINPUT1), .B(KEYINPUT94), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n326) );
  XNOR2_X1 U380 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U382 ( .A(n328), .B(n327), .Z(n338) );
  XOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT93), .Z(n330) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U386 ( .A(n332), .B(n331), .Z(n334) );
  NAND2_X1 U387 ( .A1(G225GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U391 ( .A(G155GAT), .B(G148GAT), .Z(n340) );
  XNOR2_X1 U392 ( .A(G120GAT), .B(G127GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U394 ( .A(G85GAT), .B(G162GAT), .Z(n342) );
  XNOR2_X1 U395 ( .A(G29GAT), .B(G134GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U397 ( .A(n344), .B(n343), .Z(n345) );
  XOR2_X1 U398 ( .A(n346), .B(n345), .Z(n492) );
  NOR2_X1 U399 ( .A1(n466), .A2(n492), .ZN(n447) );
  XOR2_X1 U400 ( .A(G85GAT), .B(KEYINPUT72), .Z(n385) );
  XOR2_X1 U401 ( .A(n347), .B(n385), .Z(n349) );
  NAND2_X1 U402 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n351) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n350) );
  XOR2_X1 U406 ( .A(n351), .B(n350), .Z(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n358) );
  XNOR2_X1 U408 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n354) );
  XOR2_X1 U409 ( .A(G36GAT), .B(G190GAT), .Z(n435) );
  XNOR2_X1 U410 ( .A(n354), .B(n435), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(n359), .B(G92GAT), .Z(n363) );
  XOR2_X1 U414 ( .A(G29GAT), .B(KEYINPUT7), .Z(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n366), .B(G99GAT), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n564) );
  INV_X1 U419 ( .A(KEYINPUT46), .ZN(n406) );
  XOR2_X1 U420 ( .A(KEYINPUT64), .B(KEYINPUT66), .Z(n365) );
  XNOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U423 ( .A(G1GAT), .B(G8GAT), .Z(n418) );
  XOR2_X1 U424 ( .A(n418), .B(n366), .Z(n368) );
  XNOR2_X1 U425 ( .A(G50GAT), .B(G43GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n383) );
  XOR2_X1 U428 ( .A(G22GAT), .B(G141GAT), .Z(n372) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(G197GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT67), .B(G113GAT), .Z(n374) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G15GAT), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U434 ( .A(n376), .B(n375), .Z(n381) );
  XOR2_X1 U435 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n378) );
  NAND2_X1 U436 ( .A1(G229GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U438 ( .A(KEYINPUT30), .B(n379), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n573) );
  XNOR2_X1 U441 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n384), .B(KEYINPUT13), .ZN(n410) );
  XNOR2_X1 U443 ( .A(n410), .B(n385), .ZN(n389) );
  INV_X1 U444 ( .A(n389), .ZN(n387) );
  AND2_X1 U445 ( .A1(G230GAT), .A2(G233GAT), .ZN(n388) );
  INV_X1 U446 ( .A(n388), .ZN(n386) );
  NAND2_X1 U447 ( .A1(n387), .A2(n386), .ZN(n391) );
  NAND2_X1 U448 ( .A1(n389), .A2(n388), .ZN(n390) );
  NAND2_X1 U449 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n392), .B(KEYINPUT74), .ZN(n399) );
  XOR2_X1 U451 ( .A(n393), .B(KEYINPUT32), .Z(n397) );
  XOR2_X1 U452 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n395) );
  XNOR2_X1 U453 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n394) );
  XOR2_X1 U454 ( .A(n395), .B(n394), .Z(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT73), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U456 ( .A(G204GAT), .B(G92GAT), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n439) );
  XNOR2_X1 U458 ( .A(n402), .B(n439), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n577) );
  XNOR2_X1 U460 ( .A(KEYINPUT41), .B(n577), .ZN(n553) );
  NAND2_X1 U461 ( .A1(n573), .A2(n553), .ZN(n405) );
  XOR2_X1 U462 ( .A(n406), .B(n405), .Z(n423) );
  XOR2_X1 U463 ( .A(G78GAT), .B(G211GAT), .Z(n408) );
  XNOR2_X1 U464 ( .A(G183GAT), .B(G71GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n422) );
  XOR2_X1 U466 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U467 ( .A1(G231GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U469 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n414) );
  XNOR2_X1 U470 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U472 ( .A(n416), .B(n415), .Z(n420) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U475 ( .A(n422), .B(n421), .Z(n580) );
  INV_X1 U476 ( .A(n580), .ZN(n456) );
  NAND2_X1 U477 ( .A1(n423), .A2(n456), .ZN(n424) );
  NOR2_X1 U478 ( .A1(n564), .A2(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n432) );
  XNOR2_X1 U481 ( .A(n564), .B(KEYINPUT103), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n427), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U483 ( .A1(n584), .A2(n456), .ZN(n428) );
  XNOR2_X1 U484 ( .A(KEYINPUT45), .B(n428), .ZN(n429) );
  NAND2_X1 U485 ( .A1(n429), .A2(n577), .ZN(n430) );
  NOR2_X1 U486 ( .A1(n573), .A2(n430), .ZN(n431) );
  NOR2_X1 U487 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(KEYINPUT48), .B(n433), .ZN(n528) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U490 ( .A1(G226GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT95), .Z(n441) );
  XNOR2_X1 U493 ( .A(G8GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U495 ( .A(n443), .B(n442), .Z(n495) );
  INV_X1 U496 ( .A(n495), .ZN(n521) );
  XOR2_X1 U497 ( .A(n521), .B(KEYINPUT123), .Z(n444) );
  NOR2_X1 U498 ( .A1(n528), .A2(n444), .ZN(n446) );
  AND2_X1 U499 ( .A1(n447), .A2(n570), .ZN(n450) );
  INV_X1 U500 ( .A(KEYINPUT55), .ZN(n448) );
  NOR2_X1 U501 ( .A1(n533), .A2(n451), .ZN(n565) );
  NAND2_X1 U502 ( .A1(n565), .A2(n553), .ZN(n455) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT126), .ZN(n452) );
  XNOR2_X1 U505 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n478) );
  INV_X1 U506 ( .A(n492), .ZN(n569) );
  NOR2_X1 U507 ( .A1(n564), .A2(n456), .ZN(n458) );
  XNOR2_X1 U508 ( .A(KEYINPUT16), .B(KEYINPUT78), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(n472) );
  NOR2_X1 U510 ( .A1(n533), .A2(n521), .ZN(n459) );
  NOR2_X1 U511 ( .A1(n466), .A2(n459), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT25), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(KEYINPUT96), .ZN(n464) );
  NAND2_X1 U514 ( .A1(n466), .A2(n533), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT26), .B(n462), .Z(n568) );
  XOR2_X1 U516 ( .A(n521), .B(KEYINPUT27), .Z(n467) );
  NAND2_X1 U517 ( .A1(n568), .A2(n467), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n465), .A2(n569), .ZN(n471) );
  XNOR2_X1 U520 ( .A(n466), .B(KEYINPUT28), .ZN(n503) );
  INV_X1 U521 ( .A(n503), .ZN(n531) );
  NAND2_X1 U522 ( .A1(n492), .A2(n467), .ZN(n529) );
  XOR2_X1 U523 ( .A(KEYINPUT83), .B(n498), .Z(n468) );
  NOR2_X1 U524 ( .A1(n529), .A2(n468), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n531), .A2(n469), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n488) );
  AND2_X1 U527 ( .A1(n472), .A2(n488), .ZN(n506) );
  NAND2_X1 U528 ( .A1(n577), .A2(n573), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT76), .B(n473), .Z(n490) );
  NAND2_X1 U530 ( .A1(n506), .A2(n490), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT97), .B(n474), .Z(n484) );
  NOR2_X1 U532 ( .A1(n569), .A2(n484), .ZN(n476) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U536 ( .A1(n521), .A2(n484), .ZN(n479) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n484), .A2(n533), .ZN(n483) );
  XOR2_X1 U539 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n481) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT101), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n531), .A2(n484), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(n485), .Z(n486) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NOR2_X1 U547 ( .A1(n580), .A2(n584), .ZN(n487) );
  NAND2_X1 U548 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n489), .ZN(n518) );
  NAND2_X1 U550 ( .A1(n518), .A2(n490), .ZN(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n491), .Z(n502) );
  NAND2_X1 U552 ( .A1(n492), .A2(n502), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n502), .A2(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n500) );
  NAND2_X1 U558 ( .A1(n502), .A2(n498), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n553), .ZN(n505) );
  NOR2_X1 U564 ( .A1(n573), .A2(n505), .ZN(n517) );
  NAND2_X1 U565 ( .A1(n506), .A2(n517), .ZN(n513) );
  NOR2_X1 U566 ( .A1(n569), .A2(n513), .ZN(n508) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U570 ( .A1(n521), .A2(n513), .ZN(n510) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n533), .A2(n513), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n531), .A2(n513), .ZN(n515) );
  XNOR2_X1 U576 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U580 ( .A1(n569), .A2(n525), .ZN(n520) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n533), .A2(n525), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n523), .Z(n524) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n531), .A2(n525), .ZN(n526) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n530), .B(KEYINPUT112), .ZN(n546) );
  NAND2_X1 U593 ( .A1(n531), .A2(n546), .ZN(n532) );
  NOR2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n543), .A2(n573), .ZN(n536) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT113), .Z(n534) );
  XNOR2_X1 U597 ( .A(KEYINPUT114), .B(n534), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n538) );
  NAND2_X1 U600 ( .A1(n543), .A2(n553), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n541) );
  NAND2_X1 U604 ( .A1(n543), .A2(n580), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n564), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n546), .A2(n568), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT117), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n573), .A2(n558), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT118), .B(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(n552), .Z(n555) );
  NAND2_X1 U619 ( .A1(n558), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n580), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n564), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n573), .A2(n565), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT127), .Z(n563) );
  NAND2_X1 U630 ( .A1(n565), .A2(n580), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  INV_X1 U636 ( .A(n568), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U643 ( .A(n581), .ZN(n583) );
  OR2_X1 U644 ( .A1(n583), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

