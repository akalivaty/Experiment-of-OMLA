//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT103), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G57gat), .B(G64gat), .Z(new_n205));
  AND2_X1   g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(KEYINPUT9), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n207), .B(new_n208), .Z(new_n209));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT7), .ZN(new_n211));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212));
  INV_X1    g011(.A(G85gat), .ZN(new_n213));
  INV_X1    g012(.A(G92gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(KEYINPUT8), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G99gat), .B(G106gat), .Z(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n217), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(new_n215), .A3(new_n211), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT102), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(KEYINPUT102), .A3(new_n220), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n207), .B(new_n208), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(new_n221), .A3(new_n222), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT10), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n220), .A4(new_n218), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n204), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n225), .A2(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n203), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G120gat), .B(G148gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT104), .ZN(new_n236));
  INV_X1    g035(.A(G176gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G204gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244));
  INV_X1    g043(.A(G190gat), .ZN(new_n245));
  AND2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(new_n249), .A3(new_n250), .A4(new_n245), .ZN(new_n255));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n253), .A2(new_n255), .A3(new_n256), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT70), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n262), .A2(new_n256), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n255), .A4(new_n253), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(G169gat), .B2(G176gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT65), .B(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n260), .B(new_n271), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n276), .A2(new_n245), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT24), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(G183gat), .B(G190gat), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n269), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n284));
  OAI211_X1 g083(.A(G183gat), .B(G190gat), .C1(new_n284), .C2(KEYINPUT24), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n256), .A2(KEYINPUT66), .A3(new_n279), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n276), .A2(new_n245), .A3(KEYINPUT67), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT67), .B1(new_n276), .B2(new_n245), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n260), .B1(new_n257), .B2(KEYINPUT23), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n270), .A2(G169gat), .A3(G176gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n292), .A3(KEYINPUT25), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n283), .A2(KEYINPUT68), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT68), .B1(new_n283), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n268), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297));
  OAI21_X1  g096(.A(G127gat), .B1(new_n297), .B2(KEYINPUT1), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  INV_X1    g098(.A(G127gat), .ZN(new_n300));
  INV_X1    g099(.A(G113gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G120gat), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n299), .B(new_n300), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(G134gat), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n298), .A2(G134gat), .A3(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n296), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G227gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n308), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n306), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(new_n268), .C1(new_n294), .C2(new_n295), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G15gat), .B(G43gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G71gat), .ZN(new_n319));
  INV_X1    g118(.A(G99gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n311), .B1(new_n310), .B2(new_n314), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(KEYINPUT33), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n314), .ZN(new_n327));
  INV_X1    g126(.A(new_n311), .ZN(new_n328));
  AOI221_X4 g127(.A(new_n324), .B1(KEYINPUT33), .B2(new_n321), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n317), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  INV_X1    g131(.A(new_n293), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G176gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n274), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n290), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT25), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n283), .A2(new_n293), .A3(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n313), .B1(new_n344), .B2(new_n268), .ZN(new_n345));
  INV_X1    g144(.A(new_n314), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n328), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT32), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT33), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(new_n321), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n323), .A2(new_n325), .ZN(new_n352));
  INV_X1    g151(.A(new_n316), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n315), .B(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n330), .A2(new_n331), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n352), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT74), .A3(new_n317), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n359));
  AND3_X1   g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT36), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n330), .A2(new_n362), .A3(new_n355), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(KEYINPUT72), .A3(new_n317), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT76), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(G197gat), .A2(G204gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(G197gat), .A2(G204gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT22), .ZN(new_n374));
  NAND2_X1  g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n370), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(KEYINPUT2), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n383), .A2(KEYINPUT81), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(KEYINPUT81), .ZN(new_n385));
  INV_X1    g184(.A(G148gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G141gat), .ZN(new_n387));
  INV_X1    g186(.A(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G148gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT84), .B(KEYINPUT3), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n381), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G141gat), .B(G148gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n383), .B1(new_n397), .B2(KEYINPUT82), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT83), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n380), .A2(KEYINPUT2), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n390), .B2(new_n395), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n397), .A2(KEYINPUT82), .B1(new_n380), .B2(new_n379), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n392), .B(new_n394), .C1(new_n399), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n378), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n377), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT83), .B1(new_n396), .B2(new_n398), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n403), .A3(new_n400), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n412), .A2(new_n413), .B1(new_n382), .B2(new_n391), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n407), .B(new_n409), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n408), .B(KEYINPUT87), .Z(new_n416));
  AOI21_X1  g215(.A(new_n377), .B1(new_n410), .B2(new_n405), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n376), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n376), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT88), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n368), .A3(new_n421), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n368), .A2(new_n418), .A3(new_n376), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n410), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n414), .B1(new_n424), .B2(new_n394), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n416), .B1(new_n417), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G22gat), .B(G78gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n430), .A3(new_n426), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT31), .B(G50gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G106gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n434), .A3(new_n431), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n296), .A2(new_n410), .ZN(new_n439));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n263), .B1(new_n333), .B2(new_n341), .ZN(new_n443));
  INV_X1    g242(.A(new_n440), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n442), .A3(new_n444), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n441), .A2(new_n378), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n443), .A2(new_n410), .A3(new_n440), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n296), .B2(new_n440), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n450), .A2(new_n378), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT78), .ZN(new_n454));
  INV_X1    g253(.A(G64gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(new_n214), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT30), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n452), .A2(new_n458), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n452), .A2(KEYINPUT30), .A3(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT79), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n448), .B2(new_n451), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT79), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT30), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n459), .B(new_n460), .C1(new_n462), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n392), .B1(new_n399), .B2(new_n404), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n309), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n414), .A2(new_n313), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT4), .B1(new_n469), .B2(new_n309), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n414), .A2(new_n313), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n405), .B(new_n309), .C1(new_n478), .C2(new_n414), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n467), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n313), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n474), .A2(new_n476), .B1(new_n482), .B2(new_n405), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT5), .A3(new_n467), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G57gat), .B(G85gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G1gat), .B(G29gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  INV_X1    g291(.A(new_n490), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n484), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n481), .B2(new_n484), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(KEYINPUT6), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n438), .B1(new_n466), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n244), .B1(new_n366), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n459), .ZN(new_n505));
  INV_X1    g304(.A(new_n460), .ZN(new_n506));
  AND4_X1   g305(.A1(new_n464), .A2(new_n452), .A3(KEYINPUT30), .A4(new_n458), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n464), .B1(new_n463), .B2(KEYINPUT30), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT90), .B(KEYINPUT39), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n483), .A2(new_n467), .A3(new_n510), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n470), .A2(new_n471), .A3(new_n468), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(KEYINPUT39), .C1(new_n483), .C2(new_n467), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n490), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT40), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(new_n516), .A3(new_n490), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n494), .A2(KEYINPUT91), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n481), .A2(new_n484), .A3(new_n519), .A4(new_n493), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n515), .A2(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n509), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n446), .A2(new_n447), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n444), .B1(new_n296), .B2(new_n410), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n377), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n450), .A2(new_n378), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT37), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n527), .A2(new_n457), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT92), .B(KEYINPUT37), .Z(new_n529));
  AOI21_X1  g328(.A(KEYINPUT38), .B1(new_n452), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n528), .A2(new_n530), .A3(KEYINPUT93), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT93), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n520), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n500), .B1(new_n534), .B2(new_n491), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n523), .A2(new_n524), .A3(new_n377), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n450), .A2(new_n378), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT37), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(new_n452), .ZN(new_n540));
  OAI22_X1  g339(.A1(new_n540), .A2(new_n458), .B1(KEYINPUT38), .B2(new_n463), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n522), .B(new_n438), .C1(new_n533), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n438), .ZN(new_n544));
  INV_X1    g343(.A(new_n494), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n483), .A2(new_n467), .B1(KEYINPUT5), .B2(new_n472), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT5), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n480), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n490), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n499), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n545), .B1(new_n550), .B2(new_n495), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n500), .B1(new_n551), .B2(new_n492), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n552), .B2(new_n509), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n553), .B(KEYINPUT89), .C1(new_n365), .C2(new_n360), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n504), .A2(new_n543), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n363), .A2(new_n364), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n466), .A2(new_n502), .A3(new_n556), .A4(new_n438), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n356), .A2(new_n358), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n558), .A2(new_n438), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n509), .A2(new_n535), .A3(KEYINPUT35), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT35), .A2(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n243), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT20), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT19), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n565), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G8gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(G1gat), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n570), .B1(new_n573), .B2(KEYINPUT95), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(G1gat), .B2(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI221_X1 g375(.A(new_n573), .B1(KEYINPUT95), .B2(new_n570), .C1(G1gat), .C2(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n209), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n226), .A2(KEYINPUT21), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n581), .B(new_n582), .ZN(new_n588));
  INV_X1    g387(.A(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n587), .B1(new_n585), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n569), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n588), .A2(new_n589), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n586), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n591), .A3(new_n568), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G29gat), .ZN(new_n604));
  INV_X1    g403(.A(G36gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT14), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(G29gat), .B2(G36gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT15), .ZN(new_n608));
  INV_X1    g407(.A(G43gat), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n609), .A2(G50gat), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n610), .B2(KEYINPUT94), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT14), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n607), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G43gat), .B(G50gat), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n607), .A2(new_n612), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(KEYINPUT15), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n221), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n620), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(G134gat), .ZN(new_n625));
  INV_X1    g424(.A(G134gat), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n621), .A2(new_n626), .A3(new_n622), .A4(new_n623), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n603), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n627), .A3(new_n603), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n601), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  INV_X1    g431(.A(new_n601), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n632), .A2(new_n633), .A3(new_n628), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n599), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G197gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT11), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n273), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT18), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT17), .B1(new_n616), .B2(new_n617), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n579), .B1(new_n645), .B2(KEYINPUT96), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n616), .A2(new_n617), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT96), .B1(new_n576), .B2(new_n577), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(KEYINPUT17), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G229gat), .A2(G233gat), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n653), .B(new_n643), .C1(new_n646), .C2(new_n649), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT98), .B1(new_n647), .B2(new_n579), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n647), .A2(new_n579), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n618), .A2(new_n658), .A3(new_n578), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n651), .B(KEYINPUT13), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n641), .B1(new_n655), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n650), .A2(new_n651), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n643), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n644), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n641), .A3(new_n663), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT99), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n670), .A3(new_n641), .A4(new_n663), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n664), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n636), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n563), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n502), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT105), .B(G1gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n466), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n572), .A2(new_n570), .ZN(new_n679));
  NAND2_X1  g478(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT42), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n678), .A2(new_n570), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT106), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n687));
  INV_X1    g486(.A(new_n556), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT108), .B(new_n687), .C1(new_n688), .C2(new_n361), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n360), .B2(new_n365), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n674), .A2(new_n686), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n563), .A2(new_n673), .A3(new_n558), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n686), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n674), .A2(new_n438), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n555), .A2(new_n562), .ZN(new_n702));
  INV_X1    g501(.A(new_n635), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n599), .A2(new_n672), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n704), .A2(new_n243), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n604), .A3(new_n552), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  INV_X1    g508(.A(new_n631), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n629), .A2(new_n601), .A3(new_n630), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT110), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n631), .B2(new_n634), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n543), .A2(new_n553), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n691), .B2(new_n689), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(new_n561), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n635), .B1(new_n555), .B2(new_n562), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n243), .B(KEYINPUT109), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n502), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n726), .ZN(G1328gat));
  NAND2_X1  g526(.A1(new_n707), .A2(new_n605), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n728), .A2(new_n466), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n725), .B2(new_n466), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT111), .B(KEYINPUT46), .C1(new_n728), .C2(new_n466), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(G1329gat));
  NAND2_X1  g533(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n735));
  INV_X1    g534(.A(new_n243), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n736), .A3(new_n558), .A4(new_n705), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n609), .ZN(new_n738));
  INV_X1    g537(.A(new_n692), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n735), .B(new_n738), .C1(new_n725), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n741), .B(new_n742), .Z(G1330gat));
  XOR2_X1   g542(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n544), .A3(new_n724), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n704), .A2(G50gat), .A3(new_n243), .A4(new_n706), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n544), .ZN(new_n749));
  OAI211_X1 g548(.A(KEYINPUT114), .B(new_n745), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n746), .A2(G50gat), .B1(new_n748), .B2(new_n544), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n744), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(KEYINPUT48), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(G1331gat));
  NAND2_X1  g554(.A1(new_n669), .A2(new_n671), .ZN(new_n756));
  INV_X1    g555(.A(new_n664), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n636), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n723), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT115), .Z(new_n761));
  AND2_X1   g560(.A1(new_n543), .A2(new_n553), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n561), .B1(new_n762), .B2(new_n692), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n552), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  INV_X1    g565(.A(KEYINPUT49), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n764), .B(new_n509), .C1(new_n767), .C2(new_n455), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n455), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1333gat));
  NAND3_X1  g569(.A1(new_n764), .A2(G71gat), .A3(new_n739), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n764), .A2(new_n558), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G71gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n764), .A2(new_n544), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  INV_X1    g575(.A(new_n599), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n672), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n703), .B(new_n779), .C1(new_n718), .C2(new_n561), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n692), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n778), .B1(new_n783), .B2(new_n562), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(KEYINPUT51), .A3(new_n703), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n736), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n213), .A3(new_n552), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n778), .A2(new_n736), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n722), .A2(KEYINPUT116), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT116), .B1(new_n722), .B2(new_n788), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n502), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n793), .B2(new_n213), .ZN(G1336gat));
  NAND2_X1  g593(.A1(new_n723), .A2(new_n509), .ZN(new_n795));
  AOI211_X1 g594(.A(G92gat), .B(new_n795), .C1(new_n782), .C2(new_n785), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n722), .A2(new_n788), .ZN(new_n798));
  OAI21_X1  g597(.A(G92gat), .B1(new_n798), .B2(new_n466), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n509), .B1(new_n789), .B2(new_n791), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n796), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G1337gat));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n320), .A3(new_n558), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n692), .B1(new_n790), .B2(new_n792), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n320), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(G106gat), .C1(new_n798), .C2(new_n438), .ZN(new_n809));
  INV_X1    g608(.A(new_n723), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n784), .B2(new_n703), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n763), .A2(new_n781), .A3(new_n635), .A4(new_n778), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n544), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n809), .B(new_n814), .C1(KEYINPUT117), .C2(new_n808), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n544), .B1(new_n789), .B2(new_n791), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(G106gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n818), .B2(new_n808), .ZN(G1339gat));
  NOR2_X1   g618(.A1(new_n502), .A2(new_n509), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n203), .B(new_n229), .C1(new_n232), .C2(KEYINPUT10), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n231), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n824), .B(new_n204), .C1(new_n228), .C2(new_n230), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n240), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n821), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n231), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n240), .A4(new_n825), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n241), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n672), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n656), .A2(new_n657), .A3(new_n661), .A4(new_n659), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n646), .A2(new_n649), .A3(new_n653), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n640), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT118), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n756), .A2(new_n243), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n715), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n712), .A2(new_n714), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n827), .A2(new_n241), .A3(new_n829), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n756), .A2(new_n836), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n599), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n636), .A2(new_n758), .A3(new_n243), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n820), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n559), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n672), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n846), .A2(new_n544), .A3(new_n688), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n301), .A3(new_n758), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT119), .Z(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n849), .B2(new_n810), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n303), .A3(new_n243), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  AOI21_X1  g656(.A(G127gat), .B1(new_n851), .B2(new_n599), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n777), .A2(new_n300), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n848), .B2(new_n859), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n851), .A2(new_n626), .A3(new_n703), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n635), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n559), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G134gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(G1343gat));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n544), .C1(new_n844), .C2(new_n845), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n692), .A2(new_n820), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n838), .B2(new_n831), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n837), .B(KEYINPUT121), .C1(new_n672), .C2(new_n830), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n703), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n843), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n777), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n845), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n438), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n871), .B(new_n873), .C1(new_n881), .C2(new_n870), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n882), .A2(KEYINPUT123), .A3(new_n672), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT123), .B1(new_n882), .B2(new_n672), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(G141gat), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n839), .A2(new_n843), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n845), .B1(new_n886), .B2(new_n777), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n872), .A3(new_n438), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(new_n388), .A3(new_n758), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(KEYINPUT58), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  INV_X1    g691(.A(new_n876), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n758), .A2(new_n841), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT121), .B1(new_n894), .B2(new_n837), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n635), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n599), .B1(new_n896), .B2(new_n843), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n544), .B1(new_n897), .B2(new_n845), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n872), .B1(new_n898), .B2(KEYINPUT57), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n892), .B1(new_n899), .B2(new_n871), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n758), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n889), .B1(new_n902), .B2(G141gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n891), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n386), .A3(new_n243), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n892), .A3(new_n871), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n736), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(KEYINPUT59), .A3(new_n386), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n842), .A2(new_n703), .A3(new_n841), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n599), .B1(new_n896), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n870), .B(new_n544), .C1(new_n912), .C2(new_n845), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n887), .B2(new_n438), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n913), .A2(new_n243), .A3(new_n914), .A4(new_n873), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G148gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT59), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n906), .B1(new_n910), .B2(new_n921), .ZN(G1345gat));
  AOI21_X1  g721(.A(G155gat), .B1(new_n888), .B2(new_n599), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n900), .A2(new_n901), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n777), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n924), .B2(new_n715), .ZN(new_n927));
  INV_X1    g726(.A(G162gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n739), .A2(new_n438), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n863), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT125), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n552), .A2(new_n466), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n887), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n559), .ZN(new_n936));
  OAI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n672), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n688), .A2(new_n544), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n758), .A2(new_n273), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1348gat));
  NOR3_X1   g740(.A1(new_n936), .A2(new_n337), .A3(new_n810), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n935), .A2(new_n243), .A3(new_n938), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n237), .B2(new_n943), .ZN(G1349gat));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  OAI21_X1  g744(.A(G183gat), .B1(new_n936), .B2(new_n777), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n935), .A2(new_n599), .A3(new_n254), .A4(new_n938), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n945), .A3(new_n947), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n949), .A2(KEYINPUT60), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT60), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n936), .B2(new_n635), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n840), .A2(new_n245), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n939), .B2(new_n956), .ZN(G1351gat));
  XNOR2_X1  g756(.A(KEYINPUT127), .B(G197gat), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n913), .A2(new_n914), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n692), .A3(new_n933), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n958), .B1(new_n960), .B2(new_n672), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n935), .A2(new_n929), .ZN(new_n962));
  INV_X1    g761(.A(new_n958), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(new_n758), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(G1352gat));
  NAND3_X1  g764(.A1(new_n962), .A2(new_n239), .A3(new_n243), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  OAI21_X1  g766(.A(G204gat), .B1(new_n960), .B2(new_n810), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1353gat));
  INV_X1    g768(.A(G211gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n970), .A3(new_n599), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n959), .A2(new_n599), .A3(new_n692), .A4(new_n933), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n962), .B2(new_n840), .ZN(new_n977));
  INV_X1    g776(.A(new_n960), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n703), .A2(G218gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(G1355gat));
endmodule


