

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X2 U325 ( .A(KEYINPUT48), .B(n432), .ZN(n542) );
  XNOR2_X1 U326 ( .A(KEYINPUT97), .B(n468), .ZN(n541) );
  XOR2_X1 U327 ( .A(n454), .B(n453), .Z(n526) );
  INV_X1 U328 ( .A(KEYINPUT74), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U330 ( .A(n376), .B(n375), .ZN(n377) );
  NOR2_X1 U331 ( .A1(n541), .A2(n436), .ZN(n568) );
  AND2_X1 U332 ( .A1(n455), .A2(n526), .ZN(n564) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n456) );
  XNOR2_X1 U334 ( .A(n457), .B(n456), .ZN(G1348GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n294) );
  XNOR2_X1 U336 ( .A(KEYINPUT71), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U338 ( .A(G22GAT), .B(G15GAT), .Z(n413) );
  XOR2_X1 U339 ( .A(G197GAT), .B(n413), .Z(n296) );
  XOR2_X1 U340 ( .A(G113GAT), .B(G1GAT), .Z(n341) );
  XNOR2_X1 U341 ( .A(G141GAT), .B(n341), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U343 ( .A(n298), .B(n297), .Z(n300) );
  NAND2_X1 U344 ( .A1(G229GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(n301), .B(KEYINPUT30), .Z(n304) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G8GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n302), .B(G169GAT), .ZN(n350) );
  XNOR2_X1 U349 ( .A(n350), .B(KEYINPUT68), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U351 ( .A(KEYINPUT8), .B(G50GAT), .Z(n306) );
  XNOR2_X1 U352 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(n307), .ZN(n400) );
  XNOR2_X1 U355 ( .A(n308), .B(n400), .ZN(n546) );
  INV_X1 U356 ( .A(n546), .ZN(n569) );
  XOR2_X1 U357 ( .A(n569), .B(KEYINPUT72), .Z(n529) );
  XOR2_X1 U358 ( .A(KEYINPUT3), .B(G162GAT), .Z(n310) );
  XNOR2_X1 U359 ( .A(G155GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(n311), .Z(n338) );
  XNOR2_X1 U362 ( .A(G204GAT), .B(KEYINPUT90), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n312), .B(G197GAT), .ZN(n313) );
  XOR2_X1 U364 ( .A(n313), .B(KEYINPUT21), .Z(n315) );
  XNOR2_X1 U365 ( .A(G218GAT), .B(G211GAT), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n355) );
  XOR2_X1 U367 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n317) );
  XNOR2_X1 U368 ( .A(G22GAT), .B(KEYINPUT91), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n324) );
  XOR2_X1 U370 ( .A(G106GAT), .B(G78GAT), .Z(n369) );
  XOR2_X1 U371 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n319) );
  XNOR2_X1 U372 ( .A(G148GAT), .B(G50GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n369), .B(n320), .Z(n322) );
  NAND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U377 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U378 ( .A(n355), .B(n325), .ZN(n326) );
  XOR2_X1 U379 ( .A(n338), .B(n326), .Z(n463) );
  XOR2_X1 U380 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n328) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(KEYINPUT6), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U383 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n330) );
  XNOR2_X1 U384 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U386 ( .A(n332), .B(n331), .Z(n340) );
  XOR2_X1 U387 ( .A(G127GAT), .B(KEYINPUT0), .Z(n334) );
  XNOR2_X1 U388 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n444) );
  XOR2_X1 U390 ( .A(n444), .B(KEYINPUT95), .Z(n336) );
  NAND2_X1 U391 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U395 ( .A(n342), .B(n341), .Z(n346) );
  XOR2_X1 U396 ( .A(KEYINPUT79), .B(G134GAT), .Z(n392) );
  XOR2_X1 U397 ( .A(G57GAT), .B(G120GAT), .Z(n344) );
  XNOR2_X1 U398 ( .A(G85GAT), .B(G148GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n370) );
  XNOR2_X1 U400 ( .A(n392), .B(n370), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n468) );
  XNOR2_X1 U402 ( .A(G92GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n347), .B(G176GAT), .ZN(n361) );
  XOR2_X1 U404 ( .A(KEYINPUT98), .B(n361), .Z(n349) );
  NAND2_X1 U405 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U407 ( .A(n351), .B(n350), .Z(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n353) );
  XNOR2_X1 U409 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U411 ( .A(G183GAT), .B(n354), .Z(n452) );
  XOR2_X1 U412 ( .A(n355), .B(n452), .Z(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n519) );
  INV_X1 U414 ( .A(n519), .ZN(n460) );
  XOR2_X1 U415 ( .A(n460), .B(KEYINPUT118), .Z(n433) );
  XOR2_X1 U416 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n359) );
  XNOR2_X1 U417 ( .A(KEYINPUT31), .B(KEYINPUT76), .ZN(n358) );
  XOR2_X1 U418 ( .A(n359), .B(n358), .Z(n378) );
  INV_X1 U419 ( .A(KEYINPUT32), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n363) );
  NAND2_X1 U422 ( .A1(n362), .A2(n363), .ZN(n367) );
  INV_X1 U423 ( .A(n362), .ZN(n365) );
  INV_X1 U424 ( .A(n363), .ZN(n364) );
  NAND2_X1 U425 ( .A1(n365), .A2(n364), .ZN(n366) );
  NAND2_X1 U426 ( .A1(n367), .A2(n366), .ZN(n368) );
  XOR2_X1 U427 ( .A(G99GAT), .B(G71GAT), .Z(n440) );
  XNOR2_X1 U428 ( .A(n368), .B(n440), .ZN(n372) );
  XOR2_X1 U429 ( .A(n370), .B(n369), .Z(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n417) );
  XNOR2_X1 U432 ( .A(n417), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n574) );
  XNOR2_X1 U434 ( .A(n574), .B(KEYINPUT41), .ZN(n559) );
  AND2_X1 U435 ( .A1(n546), .A2(n559), .ZN(n380) );
  XOR2_X1 U436 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n423) );
  XOR2_X1 U438 ( .A(G92GAT), .B(KEYINPUT66), .Z(n382) );
  XNOR2_X1 U439 ( .A(KEYINPUT64), .B(KEYINPUT9), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n384) );
  XNOR2_X1 U442 ( .A(G190GAT), .B(G99GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n398) );
  XOR2_X1 U445 ( .A(G106GAT), .B(KEYINPUT78), .Z(n388) );
  XNOR2_X1 U446 ( .A(G162GAT), .B(G36GAT), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n396) );
  XOR2_X1 U448 ( .A(KEYINPUT67), .B(KEYINPUT11), .Z(n390) );
  XNOR2_X1 U449 ( .A(G85GAT), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U451 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U456 ( .A(n400), .B(n399), .Z(n552) );
  XOR2_X1 U457 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n402) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(G8GAT), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n404) );
  XNOR2_X1 U461 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n421) );
  XOR2_X1 U464 ( .A(G183GAT), .B(G78GAT), .Z(n408) );
  XNOR2_X1 U465 ( .A(G155GAT), .B(G211GAT), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U467 ( .A(G64GAT), .B(G71GAT), .Z(n410) );
  XNOR2_X1 U468 ( .A(G127GAT), .B(G57GAT), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U470 ( .A(n412), .B(n411), .Z(n419) );
  XOR2_X1 U471 ( .A(KEYINPUT83), .B(n413), .Z(n415) );
  NAND2_X1 U472 ( .A1(G231GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n579) );
  INV_X1 U477 ( .A(n579), .ZN(n562) );
  OR2_X1 U478 ( .A1(n552), .A2(n562), .ZN(n422) );
  NOR2_X1 U479 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT47), .ZN(n431) );
  XOR2_X1 U481 ( .A(n552), .B(KEYINPUT104), .Z(n425) );
  XNOR2_X1 U482 ( .A(n425), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U483 ( .A1(n583), .A2(n579), .ZN(n427) );
  XNOR2_X1 U484 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  NOR2_X1 U486 ( .A1(n428), .A2(n529), .ZN(n429) );
  NAND2_X1 U487 ( .A1(n429), .A2(n574), .ZN(n430) );
  NAND2_X1 U488 ( .A1(n431), .A2(n430), .ZN(n432) );
  NAND2_X1 U489 ( .A1(n433), .A2(n542), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n434), .B(KEYINPUT54), .ZN(n435) );
  XOR2_X1 U491 ( .A(KEYINPUT119), .B(n435), .Z(n436) );
  NAND2_X1 U492 ( .A1(n463), .A2(n568), .ZN(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT55), .B(n437), .ZN(n455) );
  XOR2_X1 U494 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U495 ( .A(G113GAT), .B(G15GAT), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n443) );
  XNOR2_X1 U498 ( .A(G134GAT), .B(G43GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n448) );
  XOR2_X1 U500 ( .A(G120GAT), .B(n444), .Z(n446) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U503 ( .A(n448), .B(n447), .Z(n454) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT87), .Z(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT88), .B(G169GAT), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U508 ( .A1(n529), .A2(n564), .ZN(n457) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n480) );
  NAND2_X1 U510 ( .A1(n574), .A2(n529), .ZN(n492) );
  XOR2_X1 U511 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n459) );
  INV_X1 U512 ( .A(n552), .ZN(n537) );
  NAND2_X1 U513 ( .A1(n562), .A2(n537), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n478) );
  INV_X1 U515 ( .A(n526), .ZN(n473) );
  NOR2_X1 U516 ( .A1(n473), .A2(n460), .ZN(n461) );
  INV_X1 U517 ( .A(n463), .ZN(n470) );
  NOR2_X1 U518 ( .A1(n461), .A2(n470), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(KEYINPUT25), .ZN(n466) );
  XOR2_X1 U520 ( .A(n519), .B(KEYINPUT27), .Z(n471) );
  INV_X1 U521 ( .A(n471), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n463), .A2(n526), .ZN(n464) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(n464), .ZN(n567) );
  NAND2_X1 U524 ( .A1(n465), .A2(n567), .ZN(n543) );
  NAND2_X1 U525 ( .A1(n466), .A2(n543), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT100), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n476) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT28), .ZN(n522) );
  NOR2_X1 U529 ( .A1(n522), .A2(n471), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n472), .A2(n541), .ZN(n528) );
  XNOR2_X1 U531 ( .A(KEYINPUT99), .B(n528), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT101), .B(n477), .Z(n488) );
  NAND2_X1 U535 ( .A1(n478), .A2(n488), .ZN(n506) );
  NOR2_X1 U536 ( .A1(n492), .A2(n506), .ZN(n485) );
  NAND2_X1 U537 ( .A1(n485), .A2(n541), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n481), .Z(G1324GAT) );
  NAND2_X1 U540 ( .A1(n519), .A2(n485), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U543 ( .A1(n485), .A2(n526), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  XOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT103), .Z(n487) );
  NAND2_X1 U546 ( .A1(n485), .A2(n522), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  AND2_X1 U548 ( .A1(n579), .A2(n488), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT105), .ZN(n490) );
  NOR2_X1 U550 ( .A1(n583), .A2(n490), .ZN(n491) );
  XNOR2_X1 U551 ( .A(KEYINPUT37), .B(n491), .ZN(n516) );
  NOR2_X1 U552 ( .A1(n516), .A2(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT106), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n541), .A2(n503), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(KEYINPUT39), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n519), .A2(n503), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT108), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n501) );
  NAND2_X1 U563 ( .A1(n503), .A2(n526), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n503), .A2(n522), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(KEYINPUT110), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n569), .A2(n559), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n515), .A2(n506), .ZN(n512) );
  NAND2_X1 U572 ( .A1(n512), .A2(n541), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n519), .A2(n512), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U576 ( .A(G71GAT), .B(KEYINPUT111), .Z(n511) );
  NAND2_X1 U577 ( .A1(n512), .A2(n526), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U580 ( .A1(n512), .A2(n522), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT112), .B(n517), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n541), .A2(n523), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n519), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n526), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n542), .A2(n526), .ZN(n527) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n529), .A2(n538), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n532) );
  NAND2_X1 U598 ( .A1(n538), .A2(n559), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n535) );
  NAND2_X1 U602 ( .A1(n538), .A2(n562), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n552), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(KEYINPUT116), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n553), .A2(n546), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U614 ( .A1(n553), .A2(n559), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n562), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT117), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(n558), .Z(n561) );
  NAND2_X1 U626 ( .A1(n564), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n552), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n582), .A2(n569), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n582), .ZN(n580) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(n580), .Z(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

