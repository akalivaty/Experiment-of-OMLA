

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581;

  NOR2_X2 U320 ( .A1(n453), .A2(n565), .ZN(n439) );
  XNOR2_X1 U321 ( .A(n424), .B(n423), .ZN(n523) );
  OR2_X1 U322 ( .A1(n422), .A2(n421), .ZN(n424) );
  XNOR2_X1 U323 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n454) );
  XNOR2_X1 U324 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U325 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n341) );
  XNOR2_X1 U326 ( .A(n469), .B(n468), .ZN(n493) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n288) );
  AND2_X1 U328 ( .A1(n567), .A2(n530), .ZN(n369) );
  XNOR2_X1 U329 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U330 ( .A(KEYINPUT98), .ZN(n458) );
  XNOR2_X1 U331 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U332 ( .A(n392), .B(n288), .ZN(n356) );
  XNOR2_X1 U333 ( .A(n404), .B(n347), .ZN(n348) );
  XNOR2_X1 U334 ( .A(n356), .B(n377), .ZN(n357) );
  XNOR2_X1 U335 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U336 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U337 ( .A(n363), .B(n362), .ZN(n367) );
  XNOR2_X1 U338 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U339 ( .A(n570), .B(KEYINPUT41), .Z(n530) );
  XNOR2_X1 U340 ( .A(n543), .B(n415), .ZN(n555) );
  XOR2_X1 U341 ( .A(n435), .B(n434), .Z(n514) );
  XNOR2_X1 U342 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n474) );
  XNOR2_X1 U343 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U344 ( .A(n475), .B(n474), .ZN(G1350GAT) );
  XNOR2_X1 U345 ( .A(n473), .B(n472), .ZN(G1330GAT) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(G127GAT), .ZN(n289) );
  XNOR2_X1 U347 ( .A(n289), .B(KEYINPUT0), .ZN(n325) );
  XNOR2_X1 U348 ( .A(G120GAT), .B(G99GAT), .ZN(n290) );
  XNOR2_X1 U349 ( .A(n290), .B(G71GAT), .ZN(n364) );
  XNOR2_X1 U350 ( .A(n325), .B(n364), .ZN(n302) );
  XOR2_X1 U351 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n292) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U353 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U354 ( .A(n293), .B(G176GAT), .Z(n300) );
  XOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n295) );
  XNOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U358 ( .A(G183GAT), .B(n296), .Z(n428) );
  XOR2_X1 U359 ( .A(G169GAT), .B(G15GAT), .Z(n298) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(G43GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n346) );
  XNOR2_X1 U362 ( .A(n428), .B(n346), .ZN(n299) );
  XNOR2_X1 U363 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U364 ( .A(n302), .B(n301), .Z(n516) );
  INV_X1 U365 ( .A(n516), .ZN(n528) );
  XNOR2_X1 U366 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n303) );
  XNOR2_X1 U367 ( .A(n303), .B(KEYINPUT3), .ZN(n304) );
  XOR2_X1 U368 ( .A(n304), .B(KEYINPUT2), .Z(n306) );
  XNOR2_X1 U369 ( .A(G155GAT), .B(G162GAT), .ZN(n305) );
  XNOR2_X1 U370 ( .A(n306), .B(n305), .ZN(n326) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G22GAT), .Z(n352) );
  XOR2_X1 U372 ( .A(KEYINPUT90), .B(n352), .Z(n310) );
  XOR2_X1 U373 ( .A(G204GAT), .B(G78GAT), .Z(n308) );
  XNOR2_X1 U374 ( .A(G148GAT), .B(G106GAT), .ZN(n307) );
  XNOR2_X1 U375 ( .A(n308), .B(n307), .ZN(n365) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(n365), .ZN(n309) );
  XNOR2_X1 U377 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U378 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n312) );
  NAND2_X1 U379 ( .A1(G228GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U380 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U381 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U382 ( .A(KEYINPUT21), .B(G197GAT), .Z(n316) );
  XNOR2_X1 U383 ( .A(G218GAT), .B(KEYINPUT87), .ZN(n315) );
  XNOR2_X1 U384 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U385 ( .A(G211GAT), .B(n317), .Z(n433) );
  XNOR2_X1 U386 ( .A(n433), .B(KEYINPUT22), .ZN(n318) );
  XNOR2_X1 U387 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n326), .B(n320), .ZN(n453) );
  XOR2_X1 U389 ( .A(G113GAT), .B(G120GAT), .Z(n322) );
  XNOR2_X1 U390 ( .A(G148GAT), .B(G141GAT), .ZN(n321) );
  XNOR2_X1 U391 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U392 ( .A(G29GAT), .B(G85GAT), .Z(n323) );
  XNOR2_X1 U393 ( .A(n324), .B(n323), .ZN(n330) );
  XOR2_X1 U394 ( .A(G1GAT), .B(KEYINPUT4), .Z(n328) );
  XNOR2_X1 U395 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U396 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n330), .B(n329), .ZN(n332) );
  NAND2_X1 U398 ( .A1(G225GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n340) );
  XOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT6), .Z(n334) );
  XNOR2_X1 U401 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n333) );
  XNOR2_X1 U402 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U403 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n336) );
  XNOR2_X1 U404 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n335) );
  XNOR2_X1 U405 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U406 ( .A(n338), .B(n337), .Z(n339) );
  XOR2_X1 U407 ( .A(n340), .B(n339), .Z(n496) );
  XOR2_X1 U408 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n437) );
  XNOR2_X1 U409 ( .A(G50GAT), .B(KEYINPUT69), .ZN(n342) );
  XOR2_X1 U410 ( .A(G29GAT), .B(G36GAT), .Z(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n404) );
  XOR2_X1 U412 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n345) );
  XOR2_X1 U413 ( .A(KEYINPUT68), .B(n348), .Z(n350) );
  XOR2_X1 U414 ( .A(G1GAT), .B(G8GAT), .Z(n373) );
  XNOR2_X1 U415 ( .A(n373), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U417 ( .A(n352), .B(n351), .Z(n354) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U419 ( .A(n354), .B(n353), .Z(n567) );
  XOR2_X1 U420 ( .A(G85GAT), .B(G92GAT), .Z(n392) );
  XNOR2_X1 U421 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n355), .B(KEYINPUT71), .ZN(n377) );
  XOR2_X1 U423 ( .A(n357), .B(KEYINPUT72), .Z(n363) );
  XOR2_X1 U424 ( .A(G64GAT), .B(G176GAT), .Z(n426) );
  XNOR2_X1 U425 ( .A(n426), .B(KEYINPUT33), .ZN(n361) );
  XOR2_X1 U426 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n359) );
  XNOR2_X1 U427 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n358) );
  XNOR2_X1 U428 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n570) );
  INV_X1 U431 ( .A(KEYINPUT46), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n412) );
  XOR2_X1 U433 ( .A(G211GAT), .B(G22GAT), .Z(n371) );
  XNOR2_X1 U434 ( .A(G155GAT), .B(G78GAT), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U436 ( .A(n373), .B(n372), .Z(n375) );
  NAND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(n376), .B(KEYINPUT82), .Z(n379) );
  XNOR2_X1 U440 ( .A(n377), .B(KEYINPUT15), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U442 ( .A(G15GAT), .B(G71GAT), .Z(n381) );
  XNOR2_X1 U443 ( .A(G127GAT), .B(G183GAT), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U445 ( .A(n383), .B(n382), .Z(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n385) );
  XNOR2_X1 U447 ( .A(KEYINPUT83), .B(KEYINPUT14), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U449 ( .A(KEYINPUT84), .B(KEYINPUT80), .Z(n387) );
  XNOR2_X1 U450 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U453 ( .A(n391), .B(n390), .Z(n574) );
  XOR2_X1 U454 ( .A(G99GAT), .B(G218GAT), .Z(n394) );
  XNOR2_X1 U455 ( .A(n392), .B(KEYINPUT9), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n408) );
  XOR2_X1 U457 ( .A(G43GAT), .B(KEYINPUT10), .Z(n396) );
  XNOR2_X1 U458 ( .A(KEYINPUT11), .B(KEYINPUT67), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U460 ( .A(KEYINPUT76), .B(G190GAT), .Z(n398) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U463 ( .A(n400), .B(n399), .Z(n406) );
  XOR2_X1 U464 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n402) );
  XNOR2_X1 U465 ( .A(G162GAT), .B(G106GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U469 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U470 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XOR2_X1 U471 ( .A(n410), .B(n409), .Z(n553) );
  INV_X1 U472 ( .A(n553), .ZN(n558) );
  NOR2_X1 U473 ( .A1(n574), .A2(n558), .ZN(n411) );
  AND2_X1 U474 ( .A1(n412), .A2(n411), .ZN(n414) );
  XOR2_X1 U475 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n413) );
  XOR2_X1 U476 ( .A(n414), .B(n413), .Z(n422) );
  INV_X1 U477 ( .A(n567), .ZN(n543) );
  INV_X1 U478 ( .A(KEYINPUT70), .ZN(n415) );
  INV_X1 U479 ( .A(n570), .ZN(n444) );
  XOR2_X1 U480 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n417) );
  XOR2_X1 U481 ( .A(KEYINPUT36), .B(n553), .Z(n576) );
  NAND2_X1 U482 ( .A1(n574), .A2(n576), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n444), .A2(n418), .ZN(n419) );
  NOR2_X1 U485 ( .A1(n555), .A2(n419), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n420), .B(KEYINPUT114), .ZN(n421) );
  XNOR2_X1 U487 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n423) );
  XOR2_X1 U488 ( .A(G36GAT), .B(G92GAT), .Z(n425) );
  XOR2_X1 U489 ( .A(G169GAT), .B(G204GAT), .Z(n430) );
  NAND2_X1 U490 ( .A1(G226GAT), .A2(G233GAT), .ZN(n429) );
  XOR2_X1 U491 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n435) );
  XNOR2_X1 U493 ( .A(G8GAT), .B(n433), .ZN(n434) );
  AND2_X1 U494 ( .A1(n523), .A2(n514), .ZN(n436) );
  XOR2_X1 U495 ( .A(n437), .B(n436), .Z(n438) );
  NAND2_X1 U496 ( .A1(n496), .A2(n438), .ZN(n565) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT55), .ZN(n440) );
  NOR2_X2 U498 ( .A1(n528), .A2(n440), .ZN(n559) );
  NAND2_X1 U499 ( .A1(n559), .A2(n530), .ZN(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n441) );
  XNOR2_X1 U501 ( .A(n441), .B(G176GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(G1349GAT) );
  XOR2_X1 U503 ( .A(KEYINPUT104), .B(KEYINPUT38), .Z(n469) );
  NAND2_X1 U504 ( .A1(n444), .A2(n555), .ZN(n445) );
  XNOR2_X1 U505 ( .A(KEYINPUT75), .B(n445), .ZN(n480) );
  XOR2_X1 U506 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n467) );
  INV_X1 U507 ( .A(KEYINPUT102), .ZN(n464) );
  INV_X1 U508 ( .A(n574), .ZN(n550) );
  XOR2_X1 U509 ( .A(KEYINPUT28), .B(n453), .Z(n526) );
  INV_X1 U510 ( .A(n526), .ZN(n519) );
  XOR2_X1 U511 ( .A(n516), .B(KEYINPUT86), .Z(n446) );
  XOR2_X1 U512 ( .A(n514), .B(KEYINPUT27), .Z(n450) );
  NOR2_X1 U513 ( .A1(n496), .A2(n450), .ZN(n524) );
  NAND2_X1 U514 ( .A1(n446), .A2(n524), .ZN(n447) );
  NOR2_X1 U515 ( .A1(n519), .A2(n447), .ZN(n448) );
  XNOR2_X1 U516 ( .A(n448), .B(KEYINPUT95), .ZN(n462) );
  NAND2_X1 U517 ( .A1(n528), .A2(n453), .ZN(n449) );
  XOR2_X1 U518 ( .A(n449), .B(KEYINPUT26), .Z(n541) );
  INV_X1 U519 ( .A(n541), .ZN(n566) );
  NOR2_X1 U520 ( .A1(n566), .A2(n450), .ZN(n457) );
  INV_X1 U521 ( .A(n514), .ZN(n500) );
  NOR2_X1 U522 ( .A1(n528), .A2(n500), .ZN(n451) );
  XNOR2_X1 U523 ( .A(n451), .B(KEYINPUT96), .ZN(n452) );
  NOR2_X1 U524 ( .A1(n453), .A2(n452), .ZN(n455) );
  NOR2_X1 U525 ( .A1(n457), .A2(n456), .ZN(n459) );
  XNOR2_X1 U526 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U527 ( .A1(n460), .A2(n496), .ZN(n461) );
  NAND2_X1 U528 ( .A1(n462), .A2(n461), .ZN(n477) );
  NAND2_X1 U529 ( .A1(n550), .A2(n477), .ZN(n463) );
  XNOR2_X1 U530 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U531 ( .A1(n465), .A2(n576), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n467), .B(n466), .ZN(n510) );
  NAND2_X1 U533 ( .A1(n480), .A2(n510), .ZN(n468) );
  NAND2_X1 U534 ( .A1(n493), .A2(n516), .ZN(n473) );
  XOR2_X1 U535 ( .A(G43GAT), .B(KEYINPUT106), .Z(n471) );
  XNOR2_X1 U536 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n470) );
  NAND2_X1 U537 ( .A1(n574), .A2(n559), .ZN(n475) );
  NOR2_X1 U538 ( .A1(n558), .A2(n550), .ZN(n476) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(n476), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n479), .B(KEYINPUT99), .ZN(n495) );
  NAND2_X1 U542 ( .A1(n480), .A2(n495), .ZN(n488) );
  NOR2_X1 U543 ( .A1(n496), .A2(n488), .ZN(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U546 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  NOR2_X1 U547 ( .A1(n500), .A2(n488), .ZN(n484) );
  XOR2_X1 U548 ( .A(G8GAT), .B(n484), .Z(G1325GAT) );
  NOR2_X1 U549 ( .A1(n528), .A2(n488), .ZN(n486) );
  XNOR2_X1 U550 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U552 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  NOR2_X1 U553 ( .A1(n526), .A2(n488), .ZN(n489) );
  XOR2_X1 U554 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  INV_X1 U556 ( .A(n496), .ZN(n512) );
  NAND2_X1 U557 ( .A1(n493), .A2(n512), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n493), .A2(n514), .ZN(n492) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n493), .A2(n519), .ZN(n494) );
  XNOR2_X1 U562 ( .A(n494), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n530), .ZN(n546) );
  NOR2_X1 U564 ( .A1(n546), .A2(n567), .ZN(n509) );
  NAND2_X1 U565 ( .A1(n509), .A2(n495), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n496), .A2(n505), .ZN(n498) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n497) );
  XNOR2_X1 U568 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n500), .A2(n505), .ZN(n501) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(n501), .Z(n502) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n528), .A2(n505), .ZN(n504) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n503) );
  XNOR2_X1 U575 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n526), .A2(n505), .ZN(n507) );
  XNOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U578 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U581 ( .A(KEYINPUT111), .B(n511), .ZN(n520) );
  NAND2_X1 U582 ( .A1(n520), .A2(n512), .ZN(n513) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n514), .A2(n520), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n516), .A2(n520), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n517), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(KEYINPUT115), .B(n525), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n542), .A2(n526), .ZN(n527) );
  NOR2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n555), .A2(n537), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n532) );
  NAND2_X1 U599 ( .A1(n537), .A2(n530), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U603 ( .A1(n537), .A2(n574), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n539) );
  NAND2_X1 U607 ( .A1(n537), .A2(n558), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n552) );
  NOR2_X1 U611 ( .A1(n543), .A2(n552), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n552), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n552), .ZN(n551) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U622 ( .A1(n559), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT121), .Z(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G190GAT), .ZN(G1351GAT) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT60), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(n564), .Z(n569) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n577), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

