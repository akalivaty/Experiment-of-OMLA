

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  XOR2_X1 U322 ( .A(n448), .B(n447), .Z(n290) );
  XOR2_X1 U323 ( .A(n328), .B(n327), .Z(n291) );
  XNOR2_X1 U324 ( .A(n379), .B(KEYINPUT46), .ZN(n292) );
  XNOR2_X1 U325 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U326 ( .A(G176GAT), .B(G64GAT), .ZN(n363) );
  XNOR2_X1 U327 ( .A(n361), .B(n360), .ZN(n362) );
  NOR2_X1 U328 ( .A1(n554), .A2(n380), .ZN(n381) );
  XNOR2_X1 U329 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U330 ( .A(n373), .B(n372), .ZN(n377) );
  XNOR2_X1 U331 ( .A(n329), .B(n291), .ZN(n336) );
  XNOR2_X1 U332 ( .A(KEYINPUT102), .B(KEYINPUT36), .ZN(n340) );
  XNOR2_X1 U333 ( .A(n336), .B(n335), .ZN(n339) );
  NOR2_X1 U334 ( .A1(n526), .A2(n453), .ZN(n454) );
  XNOR2_X1 U335 ( .A(n480), .B(n340), .ZN(n580) );
  XOR2_X1 U336 ( .A(n459), .B(KEYINPUT41), .Z(n558) );
  XNOR2_X1 U337 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n458), .B(n457), .ZN(G1341GAT) );
  XNOR2_X1 U339 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n293), .B(G29GAT), .ZN(n294) );
  XOR2_X1 U341 ( .A(n294), .B(KEYINPUT7), .Z(n296) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G50GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n337) );
  XOR2_X1 U344 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n298) );
  XNOR2_X1 U345 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U347 ( .A(G113GAT), .B(G197GAT), .Z(n300) );
  XOR2_X1 U348 ( .A(G141GAT), .B(G22GAT), .Z(n435) );
  XOR2_X1 U349 ( .A(G169GAT), .B(G8GAT), .Z(n394) );
  XNOR2_X1 U350 ( .A(n435), .B(n394), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U352 ( .A(n302), .B(n301), .Z(n304) );
  NAND2_X1 U353 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U355 ( .A(n305), .B(KEYINPUT68), .Z(n308) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(G1GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n306), .B(KEYINPUT72), .ZN(n347) );
  XNOR2_X1 U358 ( .A(n347), .B(KEYINPUT29), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n337), .B(n309), .ZN(n566) );
  XNOR2_X1 U361 ( .A(KEYINPUT73), .B(n566), .ZN(n460) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n375) );
  XOR2_X1 U363 ( .A(G176GAT), .B(G190GAT), .Z(n311) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(G99GAT), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U366 ( .A(n375), .B(n312), .Z(n314) );
  NAND2_X1 U367 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U369 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n316) );
  XNOR2_X1 U370 ( .A(G169GAT), .B(G15GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U372 ( .A(n318), .B(n317), .Z(n326) );
  XOR2_X1 U373 ( .A(KEYINPUT83), .B(G134GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(G113GAT), .B(n321), .Z(n420) );
  XOR2_X1 U377 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(KEYINPUT19), .B(n324), .Z(n388) );
  XNOR2_X1 U381 ( .A(n420), .B(n388), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n476) );
  XOR2_X1 U383 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n400) );
  INV_X1 U384 ( .A(n460), .ZN(n533) );
  XOR2_X1 U385 ( .A(KEYINPUT77), .B(G162GAT), .Z(n424) );
  XOR2_X1 U386 ( .A(G190GAT), .B(G218GAT), .Z(n390) );
  XOR2_X1 U387 ( .A(n424), .B(n390), .Z(n329) );
  XOR2_X1 U388 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n328) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U390 ( .A(KEYINPUT78), .B(KEYINPUT66), .Z(n331) );
  XNOR2_X1 U391 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n334) );
  XOR2_X1 U393 ( .A(G92GAT), .B(G85GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G99GAT), .B(G106GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n367) );
  XNOR2_X1 U396 ( .A(n334), .B(n367), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n337), .B(G134GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n554) );
  XOR2_X1 U399 ( .A(KEYINPUT80), .B(n554), .Z(n480) );
  XOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT13), .Z(n374) );
  XOR2_X1 U401 ( .A(G78GAT), .B(G155GAT), .Z(n342) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U404 ( .A(n374), .B(n343), .Z(n345) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U407 ( .A(n346), .B(KEYINPUT15), .Z(n349) );
  XNOR2_X1 U408 ( .A(n347), .B(KEYINPUT12), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n357) );
  XOR2_X1 U410 ( .A(G71GAT), .B(G183GAT), .Z(n351) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G127GAT), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U413 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n353) );
  XNOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U416 ( .A(n355), .B(n354), .Z(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n536) );
  NOR2_X1 U418 ( .A1(n580), .A2(n536), .ZN(n361) );
  XNOR2_X1 U419 ( .A(KEYINPUT109), .B(KEYINPUT45), .ZN(n359) );
  INV_X1 U420 ( .A(KEYINPUT65), .ZN(n358) );
  NOR2_X1 U421 ( .A1(n533), .A2(n362), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n363), .B(KEYINPUT76), .ZN(n389) );
  XOR2_X1 U423 ( .A(G148GAT), .B(G78GAT), .Z(n423) );
  XNOR2_X1 U424 ( .A(n389), .B(n423), .ZN(n365) );
  AND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U427 ( .A(n366), .B(KEYINPUT31), .Z(n373) );
  XNOR2_X1 U428 ( .A(n367), .B(KEYINPUT33), .ZN(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n369) );
  XNOR2_X1 U430 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n368) );
  XOR2_X1 U431 ( .A(n369), .B(n368), .Z(n370) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n459) );
  NAND2_X1 U434 ( .A1(n378), .A2(n459), .ZN(n383) );
  INV_X1 U435 ( .A(n558), .ZN(n549) );
  NAND2_X1 U436 ( .A1(n566), .A2(n549), .ZN(n379) );
  NAND2_X1 U437 ( .A1(n292), .A2(n536), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(KEYINPUT47), .ZN(n382) );
  NAND2_X1 U439 ( .A1(n383), .A2(n382), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n384), .B(KEYINPUT48), .ZN(n451) );
  XOR2_X1 U441 ( .A(KEYINPUT21), .B(G211GAT), .Z(n386) );
  XNOR2_X1 U442 ( .A(KEYINPUT87), .B(G204GAT), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U444 ( .A(G197GAT), .B(n387), .ZN(n438) );
  XOR2_X1 U445 ( .A(n388), .B(n438), .Z(n398) );
  XOR2_X1 U446 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U449 ( .A(n393), .B(G92GAT), .Z(n396) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(n394), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n486) );
  NAND2_X1 U453 ( .A1(n451), .A2(n486), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n421) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n402) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(n403), .ZN(n418) );
  XOR2_X1 U459 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n405) );
  XNOR2_X1 U460 ( .A(G141GAT), .B(G120GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U462 ( .A(KEYINPUT91), .B(G57GAT), .Z(n407) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U465 ( .A(n409), .B(n408), .Z(n416) );
  XOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT3), .Z(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT88), .B(KEYINPUT2), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n427) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G162GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n427), .B(n414), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n520) );
  NAND2_X1 U476 ( .A1(n421), .A2(n520), .ZN(n422) );
  XOR2_X1 U477 ( .A(KEYINPUT64), .B(n422), .Z(n565) );
  XOR2_X1 U478 ( .A(G218GAT), .B(n423), .Z(n426) );
  XNOR2_X1 U479 ( .A(G50GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U481 ( .A(n427), .B(KEYINPUT86), .Z(n429) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U484 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n433) );
  XNOR2_X1 U486 ( .A(G106GAT), .B(KEYINPUT24), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n465) );
  NAND2_X1 U491 ( .A1(n565), .A2(n465), .ZN(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U494 ( .A1(n476), .A2(n442), .ZN(n557) );
  NOR2_X1 U495 ( .A1(n460), .A2(n557), .ZN(n444) );
  INV_X1 U496 ( .A(G169GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(G1348GAT) );
  NOR2_X1 U498 ( .A1(n536), .A2(n557), .ZN(n446) );
  INV_X1 U499 ( .A(G183GAT), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(G1350GAT) );
  NOR2_X1 U501 ( .A1(n480), .A2(n557), .ZN(n449) );
  XOR2_X1 U502 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n448) );
  XNOR2_X1 U503 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n449), .B(n290), .ZN(G1351GAT) );
  INV_X1 U505 ( .A(n476), .ZN(n526) );
  XOR2_X1 U506 ( .A(n465), .B(KEYINPUT67), .Z(n450) );
  XNOR2_X1 U507 ( .A(KEYINPUT28), .B(n450), .ZN(n530) );
  XOR2_X1 U508 ( .A(n486), .B(KEYINPUT27), .Z(n463) );
  NOR2_X1 U509 ( .A1(n463), .A2(n520), .ZN(n474) );
  NAND2_X1 U510 ( .A1(n474), .A2(n451), .ZN(n452) );
  XOR2_X1 U511 ( .A(KEYINPUT110), .B(n452), .Z(n544) );
  NAND2_X1 U512 ( .A1(n530), .A2(n544), .ZN(n453) );
  XOR2_X1 U513 ( .A(KEYINPUT111), .B(n454), .Z(n540) );
  NAND2_X1 U514 ( .A1(n540), .A2(n549), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n456) );
  XOR2_X1 U516 ( .A(G120GAT), .B(KEYINPUT113), .Z(n455) );
  INV_X1 U517 ( .A(n459), .ZN(n570) );
  NOR2_X1 U518 ( .A1(n570), .A2(n460), .ZN(n498) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n476), .A2(n465), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n543) );
  NOR2_X1 U522 ( .A1(n463), .A2(n543), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT94), .B(n464), .Z(n470) );
  NAND2_X1 U524 ( .A1(n486), .A2(n476), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT95), .ZN(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT25), .B(n468), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT96), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n472), .A2(n520), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(KEYINPUT97), .ZN(n479) );
  NAND2_X1 U532 ( .A1(n474), .A2(n530), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT92), .B(n475), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n495) );
  INV_X1 U536 ( .A(n480), .ZN(n539) );
  NOR2_X1 U537 ( .A1(n539), .A2(n536), .ZN(n481) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  NOR2_X1 U539 ( .A1(n495), .A2(n482), .ZN(n509) );
  NAND2_X1 U540 ( .A1(n498), .A2(n509), .ZN(n492) );
  NOR2_X1 U541 ( .A1(n520), .A2(n492), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  INV_X1 U545 ( .A(n486), .ZN(n523) );
  NOR2_X1 U546 ( .A1(n523), .A2(n492), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  NOR2_X1 U550 ( .A1(n526), .A2(n492), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NOR2_X1 U553 ( .A1(n530), .A2(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  NOR2_X1 U556 ( .A1(n580), .A2(n495), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n536), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n497), .ZN(n519) );
  AND2_X1 U559 ( .A1(n519), .A2(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n507) );
  NOR2_X1 U562 ( .A1(n507), .A2(n520), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n507), .A2(n523), .ZN(n504) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n507), .A2(n526), .ZN(n505) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(n505), .Z(n506) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NOR2_X1 U571 ( .A1(n507), .A2(n530), .ZN(n508) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NOR2_X1 U573 ( .A1(n558), .A2(n566), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n518), .A2(n509), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n520), .A2(n515), .ZN(n510) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n515), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n515), .ZN(n514) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n520), .A2(n529), .ZN(n521) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT106), .B(n522), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n529), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n529), .ZN(n527) );
  XOR2_X1 U594 ( .A(KEYINPUT108), .B(n527), .Z(n528) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n531), .Z(n532) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n533), .A2(n540), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  INV_X1 U602 ( .A(n536), .ZN(n573) );
  NAND2_X1 U603 ( .A1(n540), .A2(n573), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  INV_X1 U609 ( .A(n543), .ZN(n564) );
  AND2_X1 U610 ( .A1(n564), .A2(n544), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n555), .A2(n566), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U616 ( .A(KEYINPUT115), .B(n548), .Z(n551) );
  NAND2_X1 U617 ( .A1(n555), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  XOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT117), .Z(n553) );
  NAND2_X1 U620 ( .A1(n555), .A2(n573), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(KEYINPUT120), .B(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n579) );
  INV_X1 U632 ( .A(n579), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n574), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U637 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT124), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

