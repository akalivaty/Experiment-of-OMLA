//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G8gat), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  INV_X1    g006(.A(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G15gat), .ZN(new_n209));
  INV_X1    g008(.A(G15gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G22gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(G1gat), .B1(new_n209), .B2(new_n211), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n203), .B(new_n205), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n206), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n204), .A4(G8gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G64gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G57gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT93), .B(G57gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(new_n220), .ZN(new_n223));
  OR2_X1    g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT94), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT94), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n223), .A2(new_n226), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n226), .ZN(new_n233));
  INV_X1    g032(.A(G57gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G64gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n221), .A2(new_n235), .A3(KEYINPUT92), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n230), .ZN(new_n237));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT92), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n233), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n219), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT97), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n246));
  NAND2_X1  g045(.A1(G231gat), .A2(G233gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT95), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT96), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n250), .A3(new_n242), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n241), .B2(new_n242), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n248), .A3(new_n251), .ZN(new_n256));
  XNOR2_X1  g055(.A(G127gat), .B(G155gat), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n254), .B2(new_n256), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n246), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n256), .ZN(new_n261));
  INV_X1    g060(.A(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n264));
  INV_X1    g063(.A(new_n246), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G183gat), .B(G211gat), .Z(new_n267));
  AND3_X1   g066(.A1(new_n260), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n260), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n245), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n260), .A2(new_n266), .ZN(new_n271));
  INV_X1    g070(.A(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n260), .A2(new_n266), .A3(new_n267), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n244), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT98), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G99gat), .A2(G106gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT8), .ZN(new_n281));
  NAND2_X1  g080(.A1(G85gat), .A2(G92gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT7), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G85gat), .ZN(new_n285));
  INV_X1    g084(.A(G92gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n281), .A2(new_n284), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G99gat), .B(G106gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(KEYINPUT8), .A2(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n293), .A2(new_n290), .A3(new_n284), .A4(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT17), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(G36gat), .ZN(new_n299));
  INV_X1    g098(.A(G36gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT87), .ZN(new_n301));
  OAI21_X1  g100(.A(G29gat), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT14), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G29gat), .B2(G36gat), .ZN(new_n304));
  INV_X1    g103(.A(G29gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n300), .A3(KEYINPUT14), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n302), .A2(KEYINPUT15), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT15), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(KEYINPUT87), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(G36gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n304), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G43gat), .B(G50gat), .Z(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n311), .A2(new_n312), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(KEYINPUT15), .A3(new_n314), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n297), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n297), .A3(new_n318), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n296), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n296), .ZN(new_n324));
  AND2_X1   g123(.A1(G232gat), .A2(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT41), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n279), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n316), .A2(new_n297), .A3(new_n318), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n295), .B1(new_n329), .B2(new_n319), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n330), .A2(new_n278), .A3(new_n326), .A4(new_n324), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n325), .A2(KEYINPUT41), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n328), .B2(new_n331), .ZN(new_n336));
  XOR2_X1   g135(.A(G134gat), .B(G162gat), .Z(new_n337));
  NOR3_X1   g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(new_n331), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n332), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n341), .B2(new_n334), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n276), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n219), .B1(new_n329), .B2(new_n319), .ZN(new_n346));
  INV_X1    g145(.A(new_n219), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n323), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G229gat), .A2(G233gat), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n346), .A2(KEYINPUT18), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n323), .A2(new_n352), .A3(new_n347), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n219), .A2(new_n316), .A3(new_n318), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n352), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n349), .B(KEYINPUT13), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT91), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n348), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n323), .A2(new_n352), .A3(new_n347), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT91), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n357), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n351), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT18), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n348), .ZN(new_n367));
  INV_X1    g166(.A(new_n349), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n370));
  XNOR2_X1  g169(.A(G113gat), .B(G141gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT11), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G197gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT12), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n365), .B(new_n369), .C1(new_n370), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n363), .B1(new_n362), .B2(new_n357), .ZN(new_n378));
  AOI211_X1 g177(.A(KEYINPUT91), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n370), .B(new_n350), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n350), .B(new_n369), .C1(new_n378), .C2(new_n379), .ZN(new_n381));
  INV_X1    g180(.A(new_n376), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G230gat), .A2(G233gat), .ZN(new_n385));
  AND4_X1   g184(.A1(KEYINPUT99), .A2(new_n232), .A3(new_n295), .A4(new_n240), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n232), .A2(new_n240), .A3(KEYINPUT99), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT99), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n295), .B1(new_n241), .B2(new_n388), .ZN(new_n389));
  AOI211_X1 g188(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n231), .A2(new_n226), .A3(new_n229), .ZN(new_n392));
  INV_X1    g191(.A(new_n221), .ZN(new_n393));
  AND2_X1   g192(.A1(KEYINPUT93), .A2(G57gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(KEYINPUT93), .A2(G57gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n396), .B2(G64gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n227), .B1(new_n238), .B2(KEYINPUT92), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n221), .A2(new_n235), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n226), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n388), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n296), .A3(new_n387), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n398), .A2(new_n403), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT99), .A3(new_n295), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT10), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(KEYINPUT10), .A3(new_n296), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n385), .B(KEYINPUT100), .Z(new_n412));
  OAI21_X1  g211(.A(new_n391), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G120gat), .B(G148gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G176gat), .B(G204gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(KEYINPUT101), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT101), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n386), .B1(new_n389), .B2(new_n387), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n409), .B1(new_n419), .B2(KEYINPUT10), .ZN(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n390), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n416), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n385), .B1(new_n408), .B2(new_n410), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n391), .A2(new_n425), .A3(new_n423), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n417), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n384), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n345), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G57gat), .B(G85gat), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT79), .ZN(new_n431));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G120gat), .ZN(new_n437));
  INV_X1    g236(.A(G120gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G113gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G134gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G127gat), .ZN(new_n444));
  INV_X1    g243(.A(G127gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G134gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(G113gat), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n451), .A2(new_n437), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n446), .A3(new_n441), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G155gat), .B(G162gat), .Z(new_n455));
  OR2_X1    g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(KEYINPUT2), .ZN(new_n459));
  XNOR2_X1  g258(.A(G155gat), .B(G162gat), .ZN(new_n460));
  INV_X1    g259(.A(G155gat), .ZN(new_n461));
  INV_X1    g260(.A(G162gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT2), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n460), .A2(new_n456), .A3(new_n463), .A4(new_n457), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n454), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(KEYINPUT76), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT70), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n448), .B(new_n472), .C1(new_n452), .C2(new_n453), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n453), .B1(new_n437), .B2(new_n451), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n440), .A2(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT70), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT76), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n477), .A3(new_n464), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n471), .A2(new_n473), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT4), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT77), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n454), .A2(new_n465), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n474), .A2(new_n475), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(KEYINPUT3), .B2(new_n465), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT3), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n459), .A2(new_n489), .A3(new_n464), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n468), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n470), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n488), .A2(new_n490), .B1(new_n483), .B2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n479), .A2(new_n482), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n495), .A2(KEYINPUT5), .A3(new_n468), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n435), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  INV_X1    g297(.A(new_n435), .ZN(new_n499));
  INV_X1    g298(.A(new_n491), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n484), .B2(new_n485), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n498), .B(new_n499), .C1(new_n501), .C2(new_n470), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n498), .B1(new_n501), .B2(new_n470), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G64gat), .B(G92gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT74), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n515), .A2(G169gat), .A3(G176gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n516), .A2(new_n517), .B1(G169gat), .B2(G176gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(KEYINPUT66), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(G169gat), .A2(G176gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G169gat), .A2(G176gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT23), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT65), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(G183gat), .A2(G190gat), .ZN(new_n529));
  AND2_X1   g328(.A1(G183gat), .A2(G190gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(KEYINPUT24), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT64), .B1(new_n530), .B2(KEYINPUT24), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n514), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G183gat), .B2(G190gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g339(.A1(G169gat), .A2(G176gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT25), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n525), .B1(new_n519), .B2(new_n521), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G183gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT27), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT27), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G183gat), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT28), .ZN(new_n553));
  INV_X1    g352(.A(G190gat), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n523), .A2(KEYINPUT68), .A3(KEYINPUT26), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT26), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n525), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n556), .B(new_n541), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n530), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n550), .A3(new_n554), .ZN(new_n564));
  NAND2_X1  g363(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n552), .A2(new_n553), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n555), .A2(new_n562), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n513), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G197gat), .B(G204gat), .ZN(new_n572));
  INV_X1    g371(.A(G218gat), .ZN(new_n573));
  INV_X1    g372(.A(G211gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT72), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G211gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n572), .B1(new_n578), .B2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n574), .A2(G218gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n573), .A2(G211gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n573), .A2(G211gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(G218gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT73), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT22), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT72), .B(G211gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n573), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n591), .A2(new_n572), .A3(new_n586), .A4(new_n583), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n513), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n546), .B2(new_n568), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n571), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n518), .A3(new_n527), .A4(new_n524), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n544), .B1(new_n599), .B2(new_n514), .ZN(new_n600));
  INV_X1    g399(.A(new_n568), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n595), .B1(new_n602), .B2(KEYINPUT29), .ZN(new_n603));
  INV_X1    g402(.A(new_n596), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n593), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT30), .B(new_n511), .C1(new_n597), .C2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n594), .B1(new_n571), .B2(new_n596), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n604), .A3(new_n593), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n609), .A3(new_n510), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n609), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT30), .B1(new_n613), .B2(new_n511), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n507), .A2(new_n616), .A3(KEYINPUT35), .ZN(new_n617));
  XNOR2_X1  g416(.A(G78gat), .B(G106gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT31), .B(G50gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G228gat), .ZN(new_n622));
  INV_X1    g421(.A(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n588), .A2(new_n592), .A3(new_n570), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n489), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT80), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n471), .A2(new_n478), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n490), .A2(new_n570), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n593), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n626), .A2(new_n489), .B1(new_n471), .B2(new_n478), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n628), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n625), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT81), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n634), .A2(new_n628), .B1(new_n593), .B2(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n627), .A2(new_n629), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT80), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT81), .A3(new_n625), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n627), .A2(new_n465), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n632), .A2(new_n624), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n208), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  AOI211_X1 g448(.A(G22gat), .B(new_n647), .C1(new_n638), .C2(new_n643), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n621), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n476), .B(new_n473), .C1(new_n600), .C2(new_n601), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n473), .A2(new_n476), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n546), .A2(new_n653), .A3(new_n568), .ZN(new_n654));
  NAND2_X1  g453(.A1(G227gat), .A2(G233gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT71), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(KEYINPUT71), .A3(new_n658), .ZN(new_n662));
  XNOR2_X1  g461(.A(G15gat), .B(G43gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G71gat), .B(G99gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n657), .B2(KEYINPUT32), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT34), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n654), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n655), .ZN(new_n670));
  AOI211_X1 g469(.A(KEYINPUT34), .B(new_n656), .C1(new_n652), .C2(new_n654), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n657), .B(KEYINPUT32), .C1(new_n658), .C2(new_n665), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n667), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT81), .B1(new_n642), .B2(new_n625), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n637), .B(new_n624), .C1(new_n639), .C2(new_n641), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n648), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G22gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n644), .A2(new_n208), .A3(new_n648), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n681), .A3(new_n620), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n651), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n617), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT75), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n606), .A2(new_n686), .A3(new_n610), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n606), .B2(new_n610), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n614), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n504), .A2(new_n506), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT86), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n651), .A2(new_n676), .A3(new_n682), .A4(KEYINPUT86), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT35), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n685), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n690), .A2(new_n689), .B1(new_n651), .B2(new_n682), .ZN(new_n698));
  INV_X1    g497(.A(new_n675), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT36), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n667), .A2(new_n672), .A3(new_n673), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT36), .B1(new_n674), .B2(new_n675), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT82), .B1(new_n698), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n651), .A2(new_n682), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n704), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT82), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n613), .A2(new_n511), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT37), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n510), .B1(new_n613), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT37), .B1(new_n608), .B2(new_n609), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT38), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(KEYINPUT38), .A3(new_n511), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT85), .A4(KEYINPUT37), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT85), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n613), .B2(new_n712), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n507), .A2(new_n711), .A3(new_n715), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n467), .B1(new_n493), .B2(new_n494), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT39), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n499), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT83), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT83), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n727), .A3(new_n499), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n722), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(KEYINPUT39), .C1(new_n468), .C2(new_n466), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT40), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n612), .A2(new_n615), .B1(new_n435), .B2(new_n505), .ZN(new_n735));
  INV_X1    g534(.A(new_n728), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n727), .B1(new_n724), .B2(new_n499), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT40), .B(new_n731), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(KEYINPUT84), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(KEYINPUT84), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n734), .B(new_n735), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n706), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n721), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n705), .A2(new_n710), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n429), .B1(new_n697), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n507), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g546(.A1(new_n745), .A2(new_n616), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT42), .B1(new_n748), .B2(new_n202), .ZN(new_n749));
  OR2_X1    g548(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  MUX2_X1   g551(.A(KEYINPUT42), .B(new_n749), .S(new_n752), .Z(G1325gat));
  AOI21_X1  g552(.A(new_n210), .B1(new_n745), .B2(new_n704), .ZN(new_n754));
  INV_X1    g553(.A(new_n676), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(G15gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n745), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT102), .ZN(G1326gat));
  NAND2_X1  g557(.A1(new_n745), .A2(new_n706), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT43), .B(G22gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1327gat));
  AOI21_X1  g560(.A(new_n343), .B1(new_n697), .B2(new_n744), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n428), .A2(new_n276), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n305), .A3(new_n507), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n707), .A3(new_n708), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n343), .B1(new_n697), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n769), .A2(KEYINPUT44), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n617), .A2(new_n684), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n693), .A2(new_n694), .ZN(new_n772));
  INV_X1    g571(.A(new_n691), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(KEYINPUT35), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n705), .A2(new_n710), .A3(new_n743), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT44), .B(new_n344), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n763), .B(KEYINPUT103), .Z(new_n778));
  NAND3_X1  g577(.A1(new_n770), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G29gat), .B1(new_n779), .B2(new_n690), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n767), .A2(new_n780), .ZN(G1328gat));
  INV_X1    g580(.A(new_n616), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n309), .A2(new_n310), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n764), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n779), .B2(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1329gat));
  NOR3_X1   g586(.A1(new_n764), .A2(G43gat), .A3(new_n755), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n704), .A3(new_n777), .A4(new_n778), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(G43gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1330gat));
  XOR2_X1   g595(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n797));
  INV_X1    g596(.A(G50gat), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n770), .A2(new_n777), .A3(new_n778), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n706), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n742), .A2(G50gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n762), .A2(new_n763), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT107), .Z(new_n803));
  OAI21_X1  g602(.A(new_n797), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(G50gat), .B1(new_n779), .B2(new_n742), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT48), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n802), .A2(new_n807), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n805), .A2(new_n810), .A3(KEYINPUT109), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT109), .B1(new_n805), .B2(new_n810), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(G1331gat));
  NAND2_X1  g612(.A1(new_n697), .A2(new_n768), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n345), .A3(new_n384), .A4(new_n427), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT110), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n507), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(new_n222), .ZN(G1332gat));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n816), .B(new_n616), .C1(new_n819), .C2(new_n220), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n220), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(G1333gat));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n815), .B(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(G71gat), .A3(new_n755), .ZN(new_n826));
  INV_X1    g625(.A(G71gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n816), .B2(new_n704), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G71gat), .B1(new_n825), .B2(new_n708), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n816), .A2(new_n827), .A3(new_n676), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1334gat));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n706), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G78gat), .ZN(G1335gat));
  INV_X1    g634(.A(new_n276), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n377), .A2(new_n383), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n417), .A2(new_n424), .A3(new_n426), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n777), .B(new_n841), .C1(KEYINPUT44), .C2(new_n769), .ZN(new_n842));
  OAI21_X1  g641(.A(G85gat), .B1(new_n842), .B2(new_n690), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT51), .B1(new_n769), .B2(new_n838), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n507), .A2(new_n285), .A3(new_n427), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(G1336gat));
  OAI21_X1  g647(.A(G92gat), .B1(new_n842), .B2(new_n782), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n782), .A2(new_n840), .A3(G92gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n844), .B2(new_n845), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n851), .B2(KEYINPUT111), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n852), .B(new_n854), .ZN(G1337gat));
  OAI21_X1  g654(.A(G99gat), .B1(new_n842), .B2(new_n708), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n755), .A2(G99gat), .A3(new_n840), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT112), .Z(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n846), .B2(new_n858), .ZN(G1338gat));
  OAI21_X1  g658(.A(G106gat), .B1(new_n842), .B2(new_n742), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  OR3_X1    g660(.A1(new_n742), .A2(G106gat), .A3(new_n840), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n860), .B(new_n861), .C1(new_n846), .C2(new_n862), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n862), .B(KEYINPUT113), .Z(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n844), .B2(new_n845), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT114), .B1(new_n866), .B2(KEYINPUT53), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n868), .B(new_n861), .C1(new_n860), .C2(new_n865), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n863), .B1(new_n867), .B2(new_n869), .ZN(G1339gat));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n409), .B(new_n412), .C1(new_n419), .C2(KEYINPUT10), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n425), .A2(new_n873), .A3(KEYINPUT54), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n421), .B(new_n875), .C1(new_n408), .C2(new_n410), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n416), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n872), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT116), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n425), .A2(new_n873), .A3(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n416), .A3(new_n876), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n872), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n880), .A2(KEYINPUT55), .A3(new_n416), .A4(new_n876), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n426), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n837), .A2(new_n879), .A3(new_n883), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n367), .A2(new_n368), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n362), .B2(new_n357), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n375), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n365), .A2(new_n376), .A3(new_n369), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n427), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n344), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n886), .A2(new_n879), .A3(new_n883), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n891), .B(new_n890), .C1(new_n338), .C2(new_n342), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n871), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n894), .A2(new_n895), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n427), .A2(new_n890), .A3(new_n891), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n881), .A2(new_n882), .A3(new_n872), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n882), .B1(new_n881), .B2(new_n872), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(new_n885), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n902), .B2(new_n837), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT117), .B(new_n898), .C1(new_n903), .C2(new_n344), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n904), .A3(new_n276), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n345), .A2(new_n384), .A3(new_n840), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n690), .A2(new_n616), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n772), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G113gat), .B1(new_n911), .B2(new_n837), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n909), .A2(new_n683), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n384), .A2(new_n436), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1340gat));
  INV_X1    g714(.A(new_n913), .ZN(new_n916));
  OAI21_X1  g715(.A(G120gat), .B1(new_n916), .B2(new_n840), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n911), .A2(new_n449), .A3(new_n450), .A4(new_n427), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1341gat));
  OAI21_X1  g718(.A(G127gat), .B1(new_n916), .B2(new_n276), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n445), .A3(new_n836), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1342gat));
  NOR4_X1   g721(.A1(new_n276), .A2(new_n344), .A3(new_n837), .A4(new_n427), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n892), .B1(new_n894), .B2(new_n384), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n896), .B1(new_n924), .B2(new_n343), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n836), .B1(new_n925), .B2(KEYINPUT117), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n926), .B2(new_n897), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n690), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n782), .A2(new_n344), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n910), .A2(G134gat), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT118), .Z(new_n934));
  NOR2_X1   g733(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT119), .ZN(new_n936));
  OAI21_X1  g735(.A(G134gat), .B1(new_n916), .B2(new_n343), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(G1343gat));
  NOR2_X1   g737(.A1(new_n742), .A2(new_n704), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR4_X1   g739(.A1(new_n909), .A2(G141gat), .A3(new_n384), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n908), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n704), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT57), .B1(new_n907), .B2(new_n706), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n878), .A2(new_n426), .A3(new_n884), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n377), .B2(new_n383), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n343), .B1(new_n946), .B2(new_n899), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n836), .B1(new_n947), .B2(new_n898), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT57), .B(new_n706), .C1(new_n948), .C2(new_n923), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n837), .A2(new_n878), .A3(new_n886), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n344), .B1(new_n952), .B2(new_n892), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n276), .B1(new_n953), .B2(new_n896), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n742), .B1(new_n954), .B2(new_n906), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n837), .B(new_n943), .C1(new_n944), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n941), .B1(new_n958), .B2(G141gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT58), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n959), .A2(KEYINPUT121), .A3(new_n960), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT121), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(G1344gat));
  INV_X1    g763(.A(G148gat), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n944), .A2(new_n957), .ZN(new_n966));
  INV_X1    g765(.A(new_n943), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI211_X1 g767(.A(KEYINPUT59), .B(new_n965), .C1(new_n968), .C2(new_n427), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT57), .B1(new_n927), .B2(new_n742), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT57), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n971), .A2(new_n427), .A3(new_n943), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n970), .B1(new_n974), .B2(G148gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n928), .A2(new_n939), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n782), .A2(new_n965), .A3(new_n427), .ZN(new_n977));
  OAI22_X1  g776(.A1(new_n969), .A2(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G1345gat));
  NOR3_X1   g777(.A1(new_n909), .A2(new_n276), .A3(new_n940), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n979), .A2(KEYINPUT122), .ZN(new_n980));
  AOI21_X1  g779(.A(G155gat), .B1(new_n979), .B2(KEYINPUT122), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n276), .A2(new_n461), .ZN(new_n982));
  AOI22_X1  g781(.A1(new_n980), .A2(new_n981), .B1(new_n968), .B2(new_n982), .ZN(G1346gat));
  AOI21_X1  g782(.A(new_n462), .B1(new_n968), .B2(new_n344), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n976), .A2(G162gat), .A3(new_n929), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(G1347gat));
  NOR2_X1   g785(.A1(new_n507), .A2(new_n782), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n927), .A2(new_n910), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(G169gat), .B1(new_n989), .B2(new_n837), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n927), .A2(new_n683), .A3(new_n988), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n384), .A2(new_n373), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G1348gat));
  NAND3_X1  g792(.A1(new_n991), .A2(G176gat), .A3(new_n427), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT123), .ZN(new_n995));
  AOI21_X1  g794(.A(G176gat), .B1(new_n989), .B2(new_n427), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n995), .A2(new_n996), .ZN(G1349gat));
  AOI21_X1  g796(.A(new_n547), .B1(new_n991), .B2(new_n836), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n836), .A2(new_n551), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n998), .B1(new_n989), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g800(.A1(new_n989), .A2(new_n554), .A3(new_n344), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n991), .A2(new_n344), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G190gat), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n1004), .A2(KEYINPUT61), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1004), .A2(KEYINPUT61), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1351gat));
  NOR3_X1   g806(.A1(new_n927), .A2(new_n940), .A3(new_n988), .ZN(new_n1008));
  XOR2_X1   g807(.A(KEYINPUT124), .B(G197gat), .Z(new_n1009));
  NOR2_X1   g808(.A1(new_n384), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g810(.A(new_n1011), .B(KEYINPUT125), .Z(new_n1012));
  NOR2_X1   g811(.A1(new_n988), .A2(new_n704), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n742), .B1(new_n905), .B2(new_n906), .ZN(new_n1014));
  OAI211_X1 g813(.A(new_n973), .B(new_n1013), .C1(new_n1014), .C2(new_n972), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1009), .B1(new_n1015), .B2(new_n384), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1012), .A2(new_n1016), .ZN(G1352gat));
  INV_X1    g816(.A(G204gat), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1008), .A2(new_n1018), .A3(new_n427), .ZN(new_n1019));
  XOR2_X1   g818(.A(new_n1019), .B(KEYINPUT62), .Z(new_n1020));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1021));
  NOR3_X1   g820(.A1(new_n1015), .A2(new_n1021), .A3(new_n840), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1021), .B1(new_n1015), .B2(new_n840), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1023), .A2(G204gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1020), .B1(new_n1022), .B2(new_n1024), .ZN(G1353gat));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n590), .A3(new_n836), .ZN(new_n1026));
  OAI211_X1 g825(.A(KEYINPUT63), .B(G211gat), .C1(new_n1015), .C2(new_n276), .ZN(new_n1027));
  INV_X1    g826(.A(new_n1027), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n971), .A2(new_n836), .A3(new_n973), .A4(new_n1013), .ZN(new_n1029));
  AOI21_X1  g828(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1026), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1031), .A2(KEYINPUT127), .ZN(new_n1032));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1033));
  OAI211_X1 g832(.A(new_n1033), .B(new_n1026), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1032), .A2(new_n1034), .ZN(G1354gat));
  OAI21_X1  g834(.A(G218gat), .B1(new_n1015), .B2(new_n343), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n1008), .A2(new_n573), .A3(new_n344), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1036), .A2(new_n1037), .ZN(G1355gat));
endmodule


